-- Generated curve samples
-- ==================================================
-- Y_real values (no virtual zoom)
-- Curve type: sin
-- Number of samples: 2048
-- Bit range: 12 bits (0 to 4095)
-- ==================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package sin_1div4T_2048s_12b_pkg is

    type sample_array_t is array (0 to 2047) of std_logic_vector(11 downto 0);

    function vec(value : integer) return std_logic_vector;

    constant SAMPLES : sample_array_t := (
        vec(0), vec(3), vec(6), vec(9), vec(13), vec(16), vec(19), vec(22),
        vec(25), vec(28), vec(31), vec(35), vec(38), vec(41), vec(44), vec(47),
        vec(50), vec(53), vec(57), vec(60), vec(63), vec(66), vec(69), vec(72),
        vec(75), vec(79), vec(82), vec(85), vec(88), vec(91), vec(94), vec(97),
        vec(101), vec(104), vec(107), vec(110), vec(113), vec(116), vec(119), vec(123),
        vec(126), vec(129), vec(132), vec(135), vec(138), vec(141), vec(145), vec(148),
        vec(151), vec(154), vec(157), vec(160), vec(163), vec(166), vec(170), vec(173),
        vec(176), vec(179), vec(182), vec(185), vec(188), vec(192), vec(195), vec(198),
        vec(201), vec(204), vec(207), vec(210), vec(214), vec(217), vec(220), vec(223),
        vec(226), vec(229), vec(232), vec(236), vec(239), vec(242), vec(245), vec(248),
        vec(251), vec(254), vec(258), vec(261), vec(264), vec(267), vec(270), vec(273),
        vec(276), vec(279), vec(283), vec(286), vec(289), vec(292), vec(295), vec(298),
        vec(301), vec(305), vec(308), vec(311), vec(314), vec(317), vec(320), vec(323),
        vec(326), vec(330), vec(333), vec(336), vec(339), vec(342), vec(345), vec(348),
        vec(352), vec(355), vec(358), vec(361), vec(364), vec(367), vec(370), vec(373),
        vec(377), vec(380), vec(383), vec(386), vec(389), vec(392), vec(395), vec(398),
        vec(402), vec(405), vec(408), vec(411), vec(414), vec(417), vec(420), vec(423),
        vec(427), vec(430), vec(433), vec(436), vec(439), vec(442), vec(445), vec(448),
        vec(452), vec(455), vec(458), vec(461), vec(464), vec(467), vec(470), vec(473),
        vec(477), vec(480), vec(483), vec(486), vec(489), vec(492), vec(495), vec(498),
        vec(502), vec(505), vec(508), vec(511), vec(514), vec(517), vec(520), vec(523),
        vec(526), vec(530), vec(533), vec(536), vec(539), vec(542), vec(545), vec(548),
        vec(551), vec(554), vec(558), vec(561), vec(564), vec(567), vec(570), vec(573),
        vec(576), vec(579), vec(582), vec(586), vec(589), vec(592), vec(595), vec(598),
        vec(601), vec(604), vec(607), vec(610), vec(614), vec(617), vec(620), vec(623),
        vec(626), vec(629), vec(632), vec(635), vec(638), vec(642), vec(645), vec(648),
        vec(651), vec(654), vec(657), vec(660), vec(663), vec(666), vec(669), vec(673),
        vec(676), vec(679), vec(682), vec(685), vec(688), vec(691), vec(694), vec(697),
        vec(700), vec(704), vec(707), vec(710), vec(713), vec(716), vec(719), vec(722),
        vec(725), vec(728), vec(731), vec(734), vec(738), vec(741), vec(744), vec(747),
        vec(750), vec(753), vec(756), vec(759), vec(762), vec(765), vec(768), vec(772),
        vec(775), vec(778), vec(781), vec(784), vec(787), vec(790), vec(793), vec(796),
        vec(799), vec(802), vec(805), vec(809), vec(812), vec(815), vec(818), vec(821),
        vec(824), vec(827), vec(830), vec(833), vec(836), vec(839), vec(842), vec(845),
        vec(849), vec(852), vec(855), vec(858), vec(861), vec(864), vec(867), vec(870),
        vec(873), vec(876), vec(879), vec(882), vec(885), vec(888), vec(892), vec(895),
        vec(898), vec(901), vec(904), vec(907), vec(910), vec(913), vec(916), vec(919),
        vec(922), vec(925), vec(928), vec(931), vec(934), vec(937), vec(941), vec(944),
        vec(947), vec(950), vec(953), vec(956), vec(959), vec(962), vec(965), vec(968),
        vec(971), vec(974), vec(977), vec(980), vec(983), vec(986), vec(989), vec(992),
        vec(995), vec(999), vec(1002), vec(1005), vec(1008), vec(1011), vec(1014), vec(1017),
        vec(1020), vec(1023), vec(1026), vec(1029), vec(1032), vec(1035), vec(1038), vec(1041),
        vec(1044), vec(1047), vec(1050), vec(1053), vec(1056), vec(1059), vec(1062), vec(1065),
        vec(1068), vec(1071), vec(1075), vec(1078), vec(1081), vec(1084), vec(1087), vec(1090),
        vec(1093), vec(1096), vec(1099), vec(1102), vec(1105), vec(1108), vec(1111), vec(1114),
        vec(1117), vec(1120), vec(1123), vec(1126), vec(1129), vec(1132), vec(1135), vec(1138),
        vec(1141), vec(1144), vec(1147), vec(1150), vec(1153), vec(1156), vec(1159), vec(1162),
        vec(1165), vec(1168), vec(1171), vec(1174), vec(1177), vec(1180), vec(1183), vec(1186),
        vec(1189), vec(1192), vec(1195), vec(1198), vec(1201), vec(1204), vec(1207), vec(1210),
        vec(1213), vec(1216), vec(1219), vec(1222), vec(1225), vec(1228), vec(1231), vec(1234),
        vec(1237), vec(1240), vec(1243), vec(1246), vec(1249), vec(1252), vec(1255), vec(1258),
        vec(1261), vec(1264), vec(1267), vec(1270), vec(1273), vec(1276), vec(1279), vec(1282),
        vec(1285), vec(1288), vec(1291), vec(1294), vec(1297), vec(1300), vec(1303), vec(1306),
        vec(1309), vec(1312), vec(1315), vec(1318), vec(1321), vec(1324), vec(1327), vec(1330),
        vec(1333), vec(1336), vec(1339), vec(1342), vec(1345), vec(1348), vec(1351), vec(1354),
        vec(1357), vec(1359), vec(1362), vec(1365), vec(1368), vec(1371), vec(1374), vec(1377),
        vec(1380), vec(1383), vec(1386), vec(1389), vec(1392), vec(1395), vec(1398), vec(1401),
        vec(1404), vec(1407), vec(1410), vec(1413), vec(1416), vec(1419), vec(1422), vec(1424),
        vec(1427), vec(1430), vec(1433), vec(1436), vec(1439), vec(1442), vec(1445), vec(1448),
        vec(1451), vec(1454), vec(1457), vec(1460), vec(1463), vec(1466), vec(1469), vec(1472),
        vec(1474), vec(1477), vec(1480), vec(1483), vec(1486), vec(1489), vec(1492), vec(1495),
        vec(1498), vec(1501), vec(1504), vec(1507), vec(1510), vec(1512), vec(1515), vec(1518),
        vec(1521), vec(1524), vec(1527), vec(1530), vec(1533), vec(1536), vec(1539), vec(1542),
        vec(1545), vec(1547), vec(1550), vec(1553), vec(1556), vec(1559), vec(1562), vec(1565),
        vec(1568), vec(1571), vec(1574), vec(1577), vec(1579), vec(1582), vec(1585), vec(1588),
        vec(1591), vec(1594), vec(1597), vec(1600), vec(1603), vec(1605), vec(1608), vec(1611),
        vec(1614), vec(1617), vec(1620), vec(1623), vec(1626), vec(1629), vec(1631), vec(1634),
        vec(1637), vec(1640), vec(1643), vec(1646), vec(1649), vec(1652), vec(1654), vec(1657),
        vec(1660), vec(1663), vec(1666), vec(1669), vec(1672), vec(1675), vec(1677), vec(1680),
        vec(1683), vec(1686), vec(1689), vec(1692), vec(1695), vec(1697), vec(1700), vec(1703),
        vec(1706), vec(1709), vec(1712), vec(1715), vec(1717), vec(1720), vec(1723), vec(1726),
        vec(1729), vec(1732), vec(1735), vec(1737), vec(1740), vec(1743), vec(1746), vec(1749),
        vec(1752), vec(1754), vec(1757), vec(1760), vec(1763), vec(1766), vec(1769), vec(1771),
        vec(1774), vec(1777), vec(1780), vec(1783), vec(1786), vec(1788), vec(1791), vec(1794),
        vec(1797), vec(1800), vec(1803), vec(1805), vec(1808), vec(1811), vec(1814), vec(1817),
        vec(1820), vec(1822), vec(1825), vec(1828), vec(1831), vec(1834), vec(1836), vec(1839),
        vec(1842), vec(1845), vec(1848), vec(1850), vec(1853), vec(1856), vec(1859), vec(1862),
        vec(1864), vec(1867), vec(1870), vec(1873), vec(1876), vec(1878), vec(1881), vec(1884),
        vec(1887), vec(1890), vec(1892), vec(1895), vec(1898), vec(1901), vec(1903), vec(1906),
        vec(1909), vec(1912), vec(1915), vec(1917), vec(1920), vec(1923), vec(1926), vec(1928),
        vec(1931), vec(1934), vec(1937), vec(1940), vec(1942), vec(1945), vec(1948), vec(1951),
        vec(1953), vec(1956), vec(1959), vec(1962), vec(1964), vec(1967), vec(1970), vec(1973),
        vec(1975), vec(1978), vec(1981), vec(1984), vec(1986), vec(1989), vec(1992), vec(1995),
        vec(1997), vec(2000), vec(2003), vec(2006), vec(2008), vec(2011), vec(2014), vec(2017),
        vec(2019), vec(2022), vec(2025), vec(2028), vec(2030), vec(2033), vec(2036), vec(2038),
        vec(2041), vec(2044), vec(2047), vec(2049), vec(2052), vec(2055), vec(2057), vec(2060),
        vec(2063), vec(2066), vec(2068), vec(2071), vec(2074), vec(2076), vec(2079), vec(2082),
        vec(2085), vec(2087), vec(2090), vec(2093), vec(2095), vec(2098), vec(2101), vec(2103),
        vec(2106), vec(2109), vec(2112), vec(2114), vec(2117), vec(2120), vec(2122), vec(2125),
        vec(2128), vec(2130), vec(2133), vec(2136), vec(2138), vec(2141), vec(2144), vec(2146),
        vec(2149), vec(2152), vec(2154), vec(2157), vec(2160), vec(2162), vec(2165), vec(2168),
        vec(2170), vec(2173), vec(2176), vec(2178), vec(2181), vec(2184), vec(2186), vec(2189),
        vec(2192), vec(2194), vec(2197), vec(2200), vec(2202), vec(2205), vec(2208), vec(2210),
        vec(2213), vec(2216), vec(2218), vec(2221), vec(2224), vec(2226), vec(2229), vec(2231),
        vec(2234), vec(2237), vec(2239), vec(2242), vec(2245), vec(2247), vec(2250), vec(2252),
        vec(2255), vec(2258), vec(2260), vec(2263), vec(2266), vec(2268), vec(2271), vec(2273),
        vec(2276), vec(2279), vec(2281), vec(2284), vec(2286), vec(2289), vec(2292), vec(2294),
        vec(2297), vec(2299), vec(2302), vec(2305), vec(2307), vec(2310), vec(2312), vec(2315),
        vec(2318), vec(2320), vec(2323), vec(2325), vec(2328), vec(2331), vec(2333), vec(2336),
        vec(2338), vec(2341), vec(2344), vec(2346), vec(2349), vec(2351), vec(2354), vec(2356),
        vec(2359), vec(2362), vec(2364), vec(2367), vec(2369), vec(2372), vec(2374), vec(2377),
        vec(2379), vec(2382), vec(2385), vec(2387), vec(2390), vec(2392), vec(2395), vec(2397),
        vec(2400), vec(2402), vec(2405), vec(2407), vec(2410), vec(2413), vec(2415), vec(2418),
        vec(2420), vec(2423), vec(2425), vec(2428), vec(2430), vec(2433), vec(2435), vec(2438),
        vec(2440), vec(2443), vec(2445), vec(2448), vec(2450), vec(2453), vec(2456), vec(2458),
        vec(2461), vec(2463), vec(2466), vec(2468), vec(2471), vec(2473), vec(2476), vec(2478),
        vec(2481), vec(2483), vec(2486), vec(2488), vec(2491), vec(2493), vec(2496), vec(2498),
        vec(2501), vec(2503), vec(2506), vec(2508), vec(2510), vec(2513), vec(2515), vec(2518),
        vec(2520), vec(2523), vec(2525), vec(2528), vec(2530), vec(2533), vec(2535), vec(2538),
        vec(2540), vec(2543), vec(2545), vec(2548), vec(2550), vec(2552), vec(2555), vec(2557),
        vec(2560), vec(2562), vec(2565), vec(2567), vec(2570), vec(2572), vec(2575), vec(2577),
        vec(2579), vec(2582), vec(2584), vec(2587), vec(2589), vec(2592), vec(2594), vec(2596),
        vec(2599), vec(2601), vec(2604), vec(2606), vec(2609), vec(2611), vec(2613), vec(2616),
        vec(2618), vec(2621), vec(2623), vec(2626), vec(2628), vec(2630), vec(2633), vec(2635),
        vec(2638), vec(2640), vec(2642), vec(2645), vec(2647), vec(2650), vec(2652), vec(2654),
        vec(2657), vec(2659), vec(2662), vec(2664), vec(2666), vec(2669), vec(2671), vec(2673),
        vec(2676), vec(2678), vec(2681), vec(2683), vec(2685), vec(2688), vec(2690), vec(2692),
        vec(2695), vec(2697), vec(2700), vec(2702), vec(2704), vec(2707), vec(2709), vec(2711),
        vec(2714), vec(2716), vec(2718), vec(2721), vec(2723), vec(2725), vec(2728), vec(2730),
        vec(2732), vec(2735), vec(2737), vec(2739), vec(2742), vec(2744), vec(2746), vec(2749),
        vec(2751), vec(2753), vec(2756), vec(2758), vec(2760), vec(2763), vec(2765), vec(2767),
        vec(2770), vec(2772), vec(2774), vec(2777), vec(2779), vec(2781), vec(2784), vec(2786),
        vec(2788), vec(2790), vec(2793), vec(2795), vec(2797), vec(2800), vec(2802), vec(2804),
        vec(2807), vec(2809), vec(2811), vec(2813), vec(2816), vec(2818), vec(2820), vec(2822),
        vec(2825), vec(2827), vec(2829), vec(2832), vec(2834), vec(2836), vec(2838), vec(2841),
        vec(2843), vec(2845), vec(2847), vec(2850), vec(2852), vec(2854), vec(2856), vec(2859),
        vec(2861), vec(2863), vec(2865), vec(2868), vec(2870), vec(2872), vec(2874), vec(2877),
        vec(2879), vec(2881), vec(2883), vec(2886), vec(2888), vec(2890), vec(2892), vec(2894),
        vec(2897), vec(2899), vec(2901), vec(2903), vec(2906), vec(2908), vec(2910), vec(2912),
        vec(2914), vec(2917), vec(2919), vec(2921), vec(2923), vec(2925), vec(2928), vec(2930),
        vec(2932), vec(2934), vec(2936), vec(2939), vec(2941), vec(2943), vec(2945), vec(2947),
        vec(2950), vec(2952), vec(2954), vec(2956), vec(2958), vec(2960), vec(2963), vec(2965),
        vec(2967), vec(2969), vec(2971), vec(2973), vec(2976), vec(2978), vec(2980), vec(2982),
        vec(2984), vec(2986), vec(2988), vec(2991), vec(2993), vec(2995), vec(2997), vec(2999),
        vec(3001), vec(3003), vec(3006), vec(3008), vec(3010), vec(3012), vec(3014), vec(3016),
        vec(3018), vec(3021), vec(3023), vec(3025), vec(3027), vec(3029), vec(3031), vec(3033),
        vec(3035), vec(3037), vec(3040), vec(3042), vec(3044), vec(3046), vec(3048), vec(3050),
        vec(3052), vec(3054), vec(3056), vec(3058), vec(3060), vec(3063), vec(3065), vec(3067),
        vec(3069), vec(3071), vec(3073), vec(3075), vec(3077), vec(3079), vec(3081), vec(3083),
        vec(3085), vec(3087), vec(3090), vec(3092), vec(3094), vec(3096), vec(3098), vec(3100),
        vec(3102), vec(3104), vec(3106), vec(3108), vec(3110), vec(3112), vec(3114), vec(3116),
        vec(3118), vec(3120), vec(3122), vec(3124), vec(3126), vec(3128), vec(3130), vec(3132),
        vec(3134), vec(3137), vec(3139), vec(3141), vec(3143), vec(3145), vec(3147), vec(3149),
        vec(3151), vec(3153), vec(3155), vec(3157), vec(3159), vec(3161), vec(3163), vec(3165),
        vec(3167), vec(3169), vec(3171), vec(3173), vec(3175), vec(3177), vec(3179), vec(3181),
        vec(3182), vec(3184), vec(3186), vec(3188), vec(3190), vec(3192), vec(3194), vec(3196),
        vec(3198), vec(3200), vec(3202), vec(3204), vec(3206), vec(3208), vec(3210), vec(3212),
        vec(3214), vec(3216), vec(3218), vec(3220), vec(3222), vec(3224), vec(3226), vec(3227),
        vec(3229), vec(3231), vec(3233), vec(3235), vec(3237), vec(3239), vec(3241), vec(3243),
        vec(3245), vec(3247), vec(3249), vec(3251), vec(3252), vec(3254), vec(3256), vec(3258),
        vec(3260), vec(3262), vec(3264), vec(3266), vec(3268), vec(3270), vec(3271), vec(3273),
        vec(3275), vec(3277), vec(3279), vec(3281), vec(3283), vec(3285), vec(3287), vec(3288),
        vec(3290), vec(3292), vec(3294), vec(3296), vec(3298), vec(3300), vec(3301), vec(3303),
        vec(3305), vec(3307), vec(3309), vec(3311), vec(3313), vec(3314), vec(3316), vec(3318),
        vec(3320), vec(3322), vec(3324), vec(3325), vec(3327), vec(3329), vec(3331), vec(3333),
        vec(3335), vec(3336), vec(3338), vec(3340), vec(3342), vec(3344), vec(3345), vec(3347),
        vec(3349), vec(3351), vec(3353), vec(3355), vec(3356), vec(3358), vec(3360), vec(3362),
        vec(3364), vec(3365), vec(3367), vec(3369), vec(3371), vec(3372), vec(3374), vec(3376),
        vec(3378), vec(3380), vec(3381), vec(3383), vec(3385), vec(3387), vec(3388), vec(3390),
        vec(3392), vec(3394), vec(3395), vec(3397), vec(3399), vec(3401), vec(3402), vec(3404),
        vec(3406), vec(3408), vec(3409), vec(3411), vec(3413), vec(3415), vec(3416), vec(3418),
        vec(3420), vec(3422), vec(3423), vec(3425), vec(3427), vec(3428), vec(3430), vec(3432),
        vec(3434), vec(3435), vec(3437), vec(3439), vec(3440), vec(3442), vec(3444), vec(3446),
        vec(3447), vec(3449), vec(3451), vec(3452), vec(3454), vec(3456), vec(3457), vec(3459),
        vec(3461), vec(3462), vec(3464), vec(3466), vec(3467), vec(3469), vec(3471), vec(3472),
        vec(3474), vec(3476), vec(3477), vec(3479), vec(3481), vec(3482), vec(3484), vec(3486),
        vec(3487), vec(3489), vec(3491), vec(3492), vec(3494), vec(3496), vec(3497), vec(3499),
        vec(3500), vec(3502), vec(3504), vec(3505), vec(3507), vec(3509), vec(3510), vec(3512),
        vec(3513), vec(3515), vec(3517), vec(3518), vec(3520), vec(3522), vec(3523), vec(3525),
        vec(3526), vec(3528), vec(3529), vec(3531), vec(3533), vec(3534), vec(3536), vec(3537),
        vec(3539), vec(3541), vec(3542), vec(3544), vec(3545), vec(3547), vec(3548), vec(3550),
        vec(3552), vec(3553), vec(3555), vec(3556), vec(3558), vec(3559), vec(3561), vec(3562),
        vec(3564), vec(3566), vec(3567), vec(3569), vec(3570), vec(3572), vec(3573), vec(3575),
        vec(3576), vec(3578), vec(3579), vec(3581), vec(3582), vec(3584), vec(3586), vec(3587),
        vec(3589), vec(3590), vec(3592), vec(3593), vec(3595), vec(3596), vec(3598), vec(3599),
        vec(3601), vec(3602), vec(3604), vec(3605), vec(3607), vec(3608), vec(3610), vec(3611),
        vec(3612), vec(3614), vec(3615), vec(3617), vec(3618), vec(3620), vec(3621), vec(3623),
        vec(3624), vec(3626), vec(3627), vec(3629), vec(3630), vec(3632), vec(3633), vec(3634),
        vec(3636), vec(3637), vec(3639), vec(3640), vec(3642), vec(3643), vec(3645), vec(3646),
        vec(3647), vec(3649), vec(3650), vec(3652), vec(3653), vec(3655), vec(3656), vec(3657),
        vec(3659), vec(3660), vec(3662), vec(3663), vec(3664), vec(3666), vec(3667), vec(3669),
        vec(3670), vec(3671), vec(3673), vec(3674), vec(3676), vec(3677), vec(3678), vec(3680),
        vec(3681), vec(3682), vec(3684), vec(3685), vec(3687), vec(3688), vec(3689), vec(3691),
        vec(3692), vec(3693), vec(3695), vec(3696), vec(3697), vec(3699), vec(3700), vec(3701),
        vec(3703), vec(3704), vec(3705), vec(3707), vec(3708), vec(3709), vec(3711), vec(3712),
        vec(3713), vec(3715), vec(3716), vec(3717), vec(3719), vec(3720), vec(3721), vec(3723),
        vec(3724), vec(3725), vec(3727), vec(3728), vec(3729), vec(3731), vec(3732), vec(3733),
        vec(3734), vec(3736), vec(3737), vec(3738), vec(3740), vec(3741), vec(3742), vec(3743),
        vec(3745), vec(3746), vec(3747), vec(3748), vec(3750), vec(3751), vec(3752), vec(3753),
        vec(3755), vec(3756), vec(3757), vec(3758), vec(3760), vec(3761), vec(3762), vec(3763),
        vec(3765), vec(3766), vec(3767), vec(3768), vec(3770), vec(3771), vec(3772), vec(3773),
        vec(3775), vec(3776), vec(3777), vec(3778), vec(3779), vec(3781), vec(3782), vec(3783),
        vec(3784), vec(3785), vec(3787), vec(3788), vec(3789), vec(3790), vec(3791), vec(3793),
        vec(3794), vec(3795), vec(3796), vec(3797), vec(3798), vec(3800), vec(3801), vec(3802),
        vec(3803), vec(3804), vec(3805), vec(3807), vec(3808), vec(3809), vec(3810), vec(3811),
        vec(3812), vec(3814), vec(3815), vec(3816), vec(3817), vec(3818), vec(3819), vec(3820),
        vec(3821), vec(3823), vec(3824), vec(3825), vec(3826), vec(3827), vec(3828), vec(3829),
        vec(3830), vec(3832), vec(3833), vec(3834), vec(3835), vec(3836), vec(3837), vec(3838),
        vec(3839), vec(3840), vec(3841), vec(3843), vec(3844), vec(3845), vec(3846), vec(3847),
        vec(3848), vec(3849), vec(3850), vec(3851), vec(3852), vec(3853), vec(3854), vec(3855),
        vec(3856), vec(3858), vec(3859), vec(3860), vec(3861), vec(3862), vec(3863), vec(3864),
        vec(3865), vec(3866), vec(3867), vec(3868), vec(3869), vec(3870), vec(3871), vec(3872),
        vec(3873), vec(3874), vec(3875), vec(3876), vec(3877), vec(3878), vec(3879), vec(3880),
        vec(3881), vec(3882), vec(3883), vec(3884), vec(3885), vec(3886), vec(3887), vec(3888),
        vec(3889), vec(3890), vec(3891), vec(3892), vec(3893), vec(3894), vec(3895), vec(3896),
        vec(3897), vec(3898), vec(3899), vec(3900), vec(3901), vec(3902), vec(3903), vec(3904),
        vec(3905), vec(3905), vec(3906), vec(3907), vec(3908), vec(3909), vec(3910), vec(3911),
        vec(3912), vec(3913), vec(3914), vec(3915), vec(3916), vec(3917), vec(3918), vec(3918),
        vec(3919), vec(3920), vec(3921), vec(3922), vec(3923), vec(3924), vec(3925), vec(3926),
        vec(3927), vec(3928), vec(3928), vec(3929), vec(3930), vec(3931), vec(3932), vec(3933),
        vec(3934), vec(3935), vec(3935), vec(3936), vec(3937), vec(3938), vec(3939), vec(3940),
        vec(3941), vec(3941), vec(3942), vec(3943), vec(3944), vec(3945), vec(3946), vec(3947),
        vec(3947), vec(3948), vec(3949), vec(3950), vec(3951), vec(3952), vec(3952), vec(3953),
        vec(3954), vec(3955), vec(3956), vec(3956), vec(3957), vec(3958), vec(3959), vec(3960),
        vec(3960), vec(3961), vec(3962), vec(3963), vec(3964), vec(3964), vec(3965), vec(3966),
        vec(3967), vec(3968), vec(3968), vec(3969), vec(3970), vec(3971), vec(3971), vec(3972),
        vec(3973), vec(3974), vec(3974), vec(3975), vec(3976), vec(3977), vec(3977), vec(3978),
        vec(3979), vec(3980), vec(3980), vec(3981), vec(3982), vec(3983), vec(3983), vec(3984),
        vec(3985), vec(3986), vec(3986), vec(3987), vec(3988), vec(3988), vec(3989), vec(3990),
        vec(3991), vec(3991), vec(3992), vec(3993), vec(3993), vec(3994), vec(3995), vec(3995),
        vec(3996), vec(3997), vec(3997), vec(3998), vec(3999), vec(3999), vec(4000), vec(4001),
        vec(4002), vec(4002), vec(4003), vec(4003), vec(4004), vec(4005), vec(4005), vec(4006),
        vec(4007), vec(4007), vec(4008), vec(4009), vec(4009), vec(4010), vec(4011), vec(4011),
        vec(4012), vec(4013), vec(4013), vec(4014), vec(4014), vec(4015), vec(4016), vec(4016),
        vec(4017), vec(4017), vec(4018), vec(4019), vec(4019), vec(4020), vec(4020), vec(4021),
        vec(4022), vec(4022), vec(4023), vec(4023), vec(4024), vec(4025), vec(4025), vec(4026),
        vec(4026), vec(4027), vec(4027), vec(4028), vec(4029), vec(4029), vec(4030), vec(4030),
        vec(4031), vec(4031), vec(4032), vec(4032), vec(4033), vec(4034), vec(4034), vec(4035),
        vec(4035), vec(4036), vec(4036), vec(4037), vec(4037), vec(4038), vec(4038), vec(4039),
        vec(4039), vec(4040), vec(4040), vec(4041), vec(4041), vec(4042), vec(4042), vec(4043),
        vec(4043), vec(4044), vec(4044), vec(4045), vec(4045), vec(4046), vec(4046), vec(4047),
        vec(4047), vec(4048), vec(4048), vec(4049), vec(4049), vec(4050), vec(4050), vec(4051),
        vec(4051), vec(4052), vec(4052), vec(4052), vec(4053), vec(4053), vec(4054), vec(4054),
        vec(4055), vec(4055), vec(4056), vec(4056), vec(4056), vec(4057), vec(4057), vec(4058),
        vec(4058), vec(4059), vec(4059), vec(4059), vec(4060), vec(4060), vec(4061), vec(4061),
        vec(4061), vec(4062), vec(4062), vec(4063), vec(4063), vec(4063), vec(4064), vec(4064),
        vec(4065), vec(4065), vec(4065), vec(4066), vec(4066), vec(4066), vec(4067), vec(4067),
        vec(4068), vec(4068), vec(4068), vec(4069), vec(4069), vec(4069), vec(4070), vec(4070),
        vec(4070), vec(4071), vec(4071), vec(4071), vec(4072), vec(4072), vec(4072), vec(4073),
        vec(4073), vec(4073), vec(4074), vec(4074), vec(4074), vec(4075), vec(4075), vec(4075),
        vec(4076), vec(4076), vec(4076), vec(4076), vec(4077), vec(4077), vec(4077), vec(4078),
        vec(4078), vec(4078), vec(4079), vec(4079), vec(4079), vec(4079), vec(4080), vec(4080),
        vec(4080), vec(4080), vec(4081), vec(4081), vec(4081), vec(4081), vec(4082), vec(4082),
        vec(4082), vec(4082), vec(4083), vec(4083), vec(4083), vec(4083), vec(4084), vec(4084),
        vec(4084), vec(4084), vec(4085), vec(4085), vec(4085), vec(4085), vec(4085), vec(4086),
        vec(4086), vec(4086), vec(4086), vec(4086), vec(4087), vec(4087), vec(4087), vec(4087),
        vec(4087), vec(4088), vec(4088), vec(4088), vec(4088), vec(4088), vec(4089), vec(4089),
        vec(4089), vec(4089), vec(4089), vec(4089), vec(4090), vec(4090), vec(4090), vec(4090),
        vec(4090), vec(4090), vec(4091), vec(4091), vec(4091), vec(4091), vec(4091), vec(4091),
        vec(4091), vec(4091), vec(4092), vec(4092), vec(4092), vec(4092), vec(4092), vec(4092),
        vec(4092), vec(4092), vec(4093), vec(4093), vec(4093), vec(4093), vec(4093), vec(4093),
        vec(4093), vec(4093), vec(4093), vec(4093), vec(4094), vec(4094), vec(4094), vec(4094),
        vec(4094), vec(4094), vec(4094), vec(4094), vec(4094), vec(4094), vec(4094), vec(4094),
        vec(4094), vec(4094), vec(4094), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095),
        vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095),
        vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095)
    );

end package sin_1div4T_2048s_12b_pkg;

package body sin_1div4T_2048s_12b_pkg is

    function vec(value : integer) return std_logic_vector is
    begin
        return std_logic_vector(to_unsigned(value, 12));
    end function vec;

end package body sin_1div4T_2048s_12b_pkg;
