-- Generated curve samples
-- ==================================================
-- Y_real values (no virtual zoom)
-- Curve type: sin
-- Number of samples: 4096
-- Bit range: 12 bits (0 to 4095)
-- ==================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package sin_1T_4096s_12b_pkg is

    type sample_array_t is array (0 to 4095) of std_logic_vector(11 downto 0);

    function vec(value : integer) return std_logic_vector;

    constant SAMPLES : sample_array_t := (
        vec(2048), vec(2051), vec(2054), vec(2057), vec(2060), vec(2063), vec(2066), vec(2069),
        vec(2073), vec(2076), vec(2079), vec(2082), vec(2085), vec(2088), vec(2091), vec(2095),
        vec(2098), vec(2101), vec(2104), vec(2107), vec(2110), vec(2113), vec(2117), vec(2120),
        vec(2123), vec(2126), vec(2129), vec(2132), vec(2135), vec(2139), vec(2142), vec(2145),
        vec(2148), vec(2151), vec(2154), vec(2157), vec(2161), vec(2164), vec(2167), vec(2170),
        vec(2173), vec(2176), vec(2179), vec(2182), vec(2186), vec(2189), vec(2192), vec(2195),
        vec(2198), vec(2201), vec(2204), vec(2208), vec(2211), vec(2214), vec(2217), vec(2220),
        vec(2223), vec(2226), vec(2229), vec(2233), vec(2236), vec(2239), vec(2242), vec(2245),
        vec(2248), vec(2251), vec(2254), vec(2258), vec(2261), vec(2264), vec(2267), vec(2270),
        vec(2273), vec(2276), vec(2279), vec(2283), vec(2286), vec(2289), vec(2292), vec(2295),
        vec(2298), vec(2301), vec(2304), vec(2308), vec(2311), vec(2314), vec(2317), vec(2320),
        vec(2323), vec(2326), vec(2329), vec(2332), vec(2336), vec(2339), vec(2342), vec(2345),
        vec(2348), vec(2351), vec(2354), vec(2357), vec(2360), vec(2364), vec(2367), vec(2370),
        vec(2373), vec(2376), vec(2379), vec(2382), vec(2385), vec(2388), vec(2391), vec(2395),
        vec(2398), vec(2401), vec(2404), vec(2407), vec(2410), vec(2413), vec(2416), vec(2419),
        vec(2422), vec(2425), vec(2429), vec(2432), vec(2435), vec(2438), vec(2441), vec(2444),
        vec(2447), vec(2450), vec(2453), vec(2456), vec(2459), vec(2462), vec(2466), vec(2469),
        vec(2472), vec(2475), vec(2478), vec(2481), vec(2484), vec(2487), vec(2490), vec(2493),
        vec(2496), vec(2499), vec(2502), vec(2505), vec(2508), vec(2512), vec(2515), vec(2518),
        vec(2521), vec(2524), vec(2527), vec(2530), vec(2533), vec(2536), vec(2539), vec(2542),
        vec(2545), vec(2548), vec(2551), vec(2554), vec(2557), vec(2560), vec(2563), vec(2566),
        vec(2569), vec(2572), vec(2576), vec(2579), vec(2582), vec(2585), vec(2588), vec(2591),
        vec(2594), vec(2597), vec(2600), vec(2603), vec(2606), vec(2609), vec(2612), vec(2615),
        vec(2618), vec(2621), vec(2624), vec(2627), vec(2630), vec(2633), vec(2636), vec(2639),
        vec(2642), vec(2645), vec(2648), vec(2651), vec(2654), vec(2657), vec(2660), vec(2663),
        vec(2666), vec(2669), vec(2672), vec(2675), vec(2678), vec(2681), vec(2684), vec(2687),
        vec(2690), vec(2693), vec(2696), vec(2699), vec(2702), vec(2705), vec(2708), vec(2711),
        vec(2714), vec(2717), vec(2720), vec(2723), vec(2726), vec(2729), vec(2732), vec(2734),
        vec(2737), vec(2740), vec(2743), vec(2746), vec(2749), vec(2752), vec(2755), vec(2758),
        vec(2761), vec(2764), vec(2767), vec(2770), vec(2773), vec(2776), vec(2779), vec(2782),
        vec(2785), vec(2787), vec(2790), vec(2793), vec(2796), vec(2799), vec(2802), vec(2805),
        vec(2808), vec(2811), vec(2814), vec(2817), vec(2820), vec(2823), vec(2825), vec(2828),
        vec(2831), vec(2834), vec(2837), vec(2840), vec(2843), vec(2846), vec(2849), vec(2851),
        vec(2854), vec(2857), vec(2860), vec(2863), vec(2866), vec(2869), vec(2872), vec(2875),
        vec(2877), vec(2880), vec(2883), vec(2886), vec(2889), vec(2892), vec(2895), vec(2897),
        vec(2900), vec(2903), vec(2906), vec(2909), vec(2912), vec(2915), vec(2917), vec(2920),
        vec(2923), vec(2926), vec(2929), vec(2932), vec(2934), vec(2937), vec(2940), vec(2943),
        vec(2946), vec(2949), vec(2951), vec(2954), vec(2957), vec(2960), vec(2963), vec(2965),
        vec(2968), vec(2971), vec(2974), vec(2977), vec(2979), vec(2982), vec(2985), vec(2988),
        vec(2991), vec(2993), vec(2996), vec(2999), vec(3002), vec(3005), vec(3007), vec(3010),
        vec(3013), vec(3016), vec(3018), vec(3021), vec(3024), vec(3027), vec(3029), vec(3032),
        vec(3035), vec(3038), vec(3040), vec(3043), vec(3046), vec(3049), vec(3051), vec(3054),
        vec(3057), vec(3060), vec(3062), vec(3065), vec(3068), vec(3071), vec(3073), vec(3076),
        vec(3079), vec(3081), vec(3084), vec(3087), vec(3090), vec(3092), vec(3095), vec(3098),
        vec(3100), vec(3103), vec(3106), vec(3108), vec(3111), vec(3114), vec(3116), vec(3119),
        vec(3122), vec(3125), vec(3127), vec(3130), vec(3133), vec(3135), vec(3138), vec(3140),
        vec(3143), vec(3146), vec(3148), vec(3151), vec(3154), vec(3156), vec(3159), vec(3162),
        vec(3164), vec(3167), vec(3170), vec(3172), vec(3175), vec(3177), vec(3180), vec(3183),
        vec(3185), vec(3188), vec(3190), vec(3193), vec(3196), vec(3198), vec(3201), vec(3203),
        vec(3206), vec(3209), vec(3211), vec(3214), vec(3216), vec(3219), vec(3222), vec(3224),
        vec(3227), vec(3229), vec(3232), vec(3234), vec(3237), vec(3240), vec(3242), vec(3245),
        vec(3247), vec(3250), vec(3252), vec(3255), vec(3257), vec(3260), vec(3262), vec(3265),
        vec(3267), vec(3270), vec(3272), vec(3275), vec(3278), vec(3280), vec(3283), vec(3285),
        vec(3288), vec(3290), vec(3293), vec(3295), vec(3298), vec(3300), vec(3302), vec(3305),
        vec(3307), vec(3310), vec(3312), vec(3315), vec(3317), vec(3320), vec(3322), vec(3325),
        vec(3327), vec(3330), vec(3332), vec(3335), vec(3337), vec(3339), vec(3342), vec(3344),
        vec(3347), vec(3349), vec(3352), vec(3354), vec(3356), vec(3359), vec(3361), vec(3364),
        vec(3366), vec(3368), vec(3371), vec(3373), vec(3376), vec(3378), vec(3380), vec(3383),
        vec(3385), vec(3388), vec(3390), vec(3392), vec(3395), vec(3397), vec(3399), vec(3402),
        vec(3404), vec(3406), vec(3409), vec(3411), vec(3413), vec(3416), vec(3418), vec(3420),
        vec(3423), vec(3425), vec(3427), vec(3430), vec(3432), vec(3434), vec(3437), vec(3439),
        vec(3441), vec(3444), vec(3446), vec(3448), vec(3450), vec(3453), vec(3455), vec(3457),
        vec(3460), vec(3462), vec(3464), vec(3466), vec(3469), vec(3471), vec(3473), vec(3475),
        vec(3478), vec(3480), vec(3482), vec(3484), vec(3487), vec(3489), vec(3491), vec(3493),
        vec(3496), vec(3498), vec(3500), vec(3502), vec(3504), vec(3507), vec(3509), vec(3511),
        vec(3513), vec(3515), vec(3518), vec(3520), vec(3522), vec(3524), vec(3526), vec(3529),
        vec(3531), vec(3533), vec(3535), vec(3537), vec(3539), vec(3541), vec(3544), vec(3546),
        vec(3548), vec(3550), vec(3552), vec(3554), vec(3556), vec(3559), vec(3561), vec(3563),
        vec(3565), vec(3567), vec(3569), vec(3571), vec(3573), vec(3575), vec(3577), vec(3580),
        vec(3582), vec(3584), vec(3586), vec(3588), vec(3590), vec(3592), vec(3594), vec(3596),
        vec(3598), vec(3600), vec(3602), vec(3604), vec(3606), vec(3608), vec(3610), vec(3612),
        vec(3614), vec(3616), vec(3618), vec(3621), vec(3623), vec(3625), vec(3627), vec(3629),
        vec(3631), vec(3633), vec(3634), vec(3636), vec(3638), vec(3640), vec(3642), vec(3644),
        vec(3646), vec(3648), vec(3650), vec(3652), vec(3654), vec(3656), vec(3658), vec(3660),
        vec(3662), vec(3664), vec(3666), vec(3668), vec(3670), vec(3672), vec(3673), vec(3675),
        vec(3677), vec(3679), vec(3681), vec(3683), vec(3685), vec(3687), vec(3689), vec(3690),
        vec(3692), vec(3694), vec(3696), vec(3698), vec(3700), vec(3702), vec(3704), vec(3705),
        vec(3707), vec(3709), vec(3711), vec(3713), vec(3715), vec(3716), vec(3718), vec(3720),
        vec(3722), vec(3724), vec(3725), vec(3727), vec(3729), vec(3731), vec(3733), vec(3734),
        vec(3736), vec(3738), vec(3740), vec(3741), vec(3743), vec(3745), vec(3747), vec(3748),
        vec(3750), vec(3752), vec(3754), vec(3755), vec(3757), vec(3759), vec(3761), vec(3762),
        vec(3764), vec(3766), vec(3767), vec(3769), vec(3771), vec(3773), vec(3774), vec(3776),
        vec(3778), vec(3779), vec(3781), vec(3783), vec(3784), vec(3786), vec(3788), vec(3789),
        vec(3791), vec(3793), vec(3794), vec(3796), vec(3797), vec(3799), vec(3801), vec(3802),
        vec(3804), vec(3806), vec(3807), vec(3809), vec(3810), vec(3812), vec(3814), vec(3815),
        vec(3817), vec(3818), vec(3820), vec(3821), vec(3823), vec(3825), vec(3826), vec(3828),
        vec(3829), vec(3831), vec(3832), vec(3834), vec(3835), vec(3837), vec(3838), vec(3840),
        vec(3842), vec(3843), vec(3845), vec(3846), vec(3848), vec(3849), vec(3851), vec(3852),
        vec(3853), vec(3855), vec(3856), vec(3858), vec(3859), vec(3861), vec(3862), vec(3864),
        vec(3865), vec(3867), vec(3868), vec(3870), vec(3871), vec(3872), vec(3874), vec(3875),
        vec(3877), vec(3878), vec(3879), vec(3881), vec(3882), vec(3884), vec(3885), vec(3886),
        vec(3888), vec(3889), vec(3891), vec(3892), vec(3893), vec(3895), vec(3896), vec(3897),
        vec(3899), vec(3900), vec(3901), vec(3903), vec(3904), vec(3905), vec(3907), vec(3908),
        vec(3909), vec(3911), vec(3912), vec(3913), vec(3914), vec(3916), vec(3917), vec(3918),
        vec(3920), vec(3921), vec(3922), vec(3923), vec(3925), vec(3926), vec(3927), vec(3928),
        vec(3930), vec(3931), vec(3932), vec(3933), vec(3935), vec(3936), vec(3937), vec(3938),
        vec(3939), vec(3941), vec(3942), vec(3943), vec(3944), vec(3945), vec(3946), vec(3948),
        vec(3949), vec(3950), vec(3951), vec(3952), vec(3953), vec(3955), vec(3956), vec(3957),
        vec(3958), vec(3959), vec(3960), vec(3961), vec(3963), vec(3964), vec(3965), vec(3966),
        vec(3967), vec(3968), vec(3969), vec(3970), vec(3971), vec(3972), vec(3973), vec(3974),
        vec(3976), vec(3977), vec(3978), vec(3979), vec(3980), vec(3981), vec(3982), vec(3983),
        vec(3984), vec(3985), vec(3986), vec(3987), vec(3988), vec(3989), vec(3990), vec(3991),
        vec(3992), vec(3993), vec(3994), vec(3995), vec(3996), vec(3997), vec(3998), vec(3999),
        vec(4000), vec(4001), vec(4001), vec(4002), vec(4003), vec(4004), vec(4005), vec(4006),
        vec(4007), vec(4008), vec(4009), vec(4010), vec(4011), vec(4012), vec(4012), vec(4013),
        vec(4014), vec(4015), vec(4016), vec(4017), vec(4018), vec(4018), vec(4019), vec(4020),
        vec(4021), vec(4022), vec(4023), vec(4023), vec(4024), vec(4025), vec(4026), vec(4027),
        vec(4028), vec(4028), vec(4029), vec(4030), vec(4031), vec(4031), vec(4032), vec(4033),
        vec(4034), vec(4035), vec(4035), vec(4036), vec(4037), vec(4038), vec(4038), vec(4039),
        vec(4040), vec(4040), vec(4041), vec(4042), vec(4043), vec(4043), vec(4044), vec(4045),
        vec(4045), vec(4046), vec(4047), vec(4047), vec(4048), vec(4049), vec(4049), vec(4050),
        vec(4051), vec(4051), vec(4052), vec(4053), vec(4053), vec(4054), vec(4055), vec(4055),
        vec(4056), vec(4056), vec(4057), vec(4058), vec(4058), vec(4059), vec(4059), vec(4060),
        vec(4061), vec(4061), vec(4062), vec(4062), vec(4063), vec(4063), vec(4064), vec(4064),
        vec(4065), vec(4066), vec(4066), vec(4067), vec(4067), vec(4068), vec(4068), vec(4069),
        vec(4069), vec(4070), vec(4070), vec(4071), vec(4071), vec(4072), vec(4072), vec(4072),
        vec(4073), vec(4073), vec(4074), vec(4074), vec(4075), vec(4075), vec(4076), vec(4076),
        vec(4076), vec(4077), vec(4077), vec(4078), vec(4078), vec(4079), vec(4079), vec(4079),
        vec(4080), vec(4080), vec(4080), vec(4081), vec(4081), vec(4082), vec(4082), vec(4082),
        vec(4083), vec(4083), vec(4083), vec(4084), vec(4084), vec(4084), vec(4085), vec(4085),
        vec(4085), vec(4086), vec(4086), vec(4086), vec(4086), vec(4087), vec(4087), vec(4087),
        vec(4088), vec(4088), vec(4088), vec(4088), vec(4089), vec(4089), vec(4089), vec(4089),
        vec(4090), vec(4090), vec(4090), vec(4090), vec(4090), vec(4091), vec(4091), vec(4091),
        vec(4091), vec(4091), vec(4092), vec(4092), vec(4092), vec(4092), vec(4092), vec(4092),
        vec(4093), vec(4093), vec(4093), vec(4093), vec(4093), vec(4093), vec(4093), vec(4094),
        vec(4094), vec(4094), vec(4094), vec(4094), vec(4094), vec(4094), vec(4094), vec(4094),
        vec(4094), vec(4094), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095),
        vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095),
        vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095),
        vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4094),
        vec(4094), vec(4094), vec(4094), vec(4094), vec(4094), vec(4094), vec(4094), vec(4094),
        vec(4094), vec(4093), vec(4093), vec(4093), vec(4093), vec(4093), vec(4093), vec(4093),
        vec(4092), vec(4092), vec(4092), vec(4092), vec(4092), vec(4092), vec(4091), vec(4091),
        vec(4091), vec(4091), vec(4091), vec(4090), vec(4090), vec(4090), vec(4090), vec(4090),
        vec(4089), vec(4089), vec(4089), vec(4089), vec(4088), vec(4088), vec(4088), vec(4088),
        vec(4087), vec(4087), vec(4087), vec(4087), vec(4086), vec(4086), vec(4086), vec(4085),
        vec(4085), vec(4085), vec(4084), vec(4084), vec(4084), vec(4083), vec(4083), vec(4083),
        vec(4082), vec(4082), vec(4082), vec(4081), vec(4081), vec(4081), vec(4080), vec(4080),
        vec(4079), vec(4079), vec(4079), vec(4078), vec(4078), vec(4078), vec(4077), vec(4077),
        vec(4076), vec(4076), vec(4075), vec(4075), vec(4075), vec(4074), vec(4074), vec(4073),
        vec(4073), vec(4072), vec(4072), vec(4071), vec(4071), vec(4070), vec(4070), vec(4069),
        vec(4069), vec(4068), vec(4068), vec(4067), vec(4067), vec(4066), vec(4066), vec(4065),
        vec(4065), vec(4064), vec(4064), vec(4063), vec(4063), vec(4062), vec(4061), vec(4061),
        vec(4060), vec(4060), vec(4059), vec(4058), vec(4058), vec(4057), vec(4057), vec(4056),
        vec(4055), vec(4055), vec(4054), vec(4054), vec(4053), vec(4052), vec(4052), vec(4051),
        vec(4050), vec(4050), vec(4049), vec(4048), vec(4048), vec(4047), vec(4046), vec(4046),
        vec(4045), vec(4044), vec(4044), vec(4043), vec(4042), vec(4042), vec(4041), vec(4040),
        vec(4039), vec(4039), vec(4038), vec(4037), vec(4036), vec(4036), vec(4035), vec(4034),
        vec(4033), vec(4033), vec(4032), vec(4031), vec(4030), vec(4030), vec(4029), vec(4028),
        vec(4027), vec(4026), vec(4026), vec(4025), vec(4024), vec(4023), vec(4022), vec(4021),
        vec(4021), vec(4020), vec(4019), vec(4018), vec(4017), vec(4016), vec(4015), vec(4015),
        vec(4014), vec(4013), vec(4012), vec(4011), vec(4010), vec(4009), vec(4008), vec(4007),
        vec(4007), vec(4006), vec(4005), vec(4004), vec(4003), vec(4002), vec(4001), vec(4000),
        vec(3999), vec(3998), vec(3997), vec(3996), vec(3995), vec(3994), vec(3993), vec(3992),
        vec(3991), vec(3990), vec(3989), vec(3988), vec(3987), vec(3986), vec(3985), vec(3984),
        vec(3983), vec(3982), vec(3981), vec(3980), vec(3979), vec(3978), vec(3977), vec(3976),
        vec(3975), vec(3974), vec(3973), vec(3972), vec(3971), vec(3970), vec(3969), vec(3967),
        vec(3966), vec(3965), vec(3964), vec(3963), vec(3962), vec(3961), vec(3960), vec(3959),
        vec(3957), vec(3956), vec(3955), vec(3954), vec(3953), vec(3952), vec(3951), vec(3949),
        vec(3948), vec(3947), vec(3946), vec(3945), vec(3944), vec(3942), vec(3941), vec(3940),
        vec(3939), vec(3938), vec(3936), vec(3935), vec(3934), vec(3933), vec(3931), vec(3930),
        vec(3929), vec(3928), vec(3927), vec(3925), vec(3924), vec(3923), vec(3921), vec(3920),
        vec(3919), vec(3918), vec(3916), vec(3915), vec(3914), vec(3913), vec(3911), vec(3910),
        vec(3909), vec(3907), vec(3906), vec(3905), vec(3903), vec(3902), vec(3901), vec(3899),
        vec(3898), vec(3897), vec(3895), vec(3894), vec(3893), vec(3891), vec(3890), vec(3888),
        vec(3887), vec(3886), vec(3884), vec(3883), vec(3882), vec(3880), vec(3879), vec(3877),
        vec(3876), vec(3875), vec(3873), vec(3872), vec(3870), vec(3869), vec(3867), vec(3866),
        vec(3864), vec(3863), vec(3862), vec(3860), vec(3859), vec(3857), vec(3856), vec(3854),
        vec(3853), vec(3851), vec(3850), vec(3848), vec(3847), vec(3845), vec(3844), vec(3842),
        vec(3841), vec(3839), vec(3838), vec(3836), vec(3835), vec(3833), vec(3832), vec(3830),
        vec(3828), vec(3827), vec(3825), vec(3824), vec(3822), vec(3821), vec(3819), vec(3818),
        vec(3816), vec(3814), vec(3813), vec(3811), vec(3810), vec(3808), vec(3806), vec(3805),
        vec(3803), vec(3802), vec(3800), vec(3798), vec(3797), vec(3795), vec(3793), vec(3792),
        vec(3790), vec(3788), vec(3787), vec(3785), vec(3783), vec(3782), vec(3780), vec(3778),
        vec(3777), vec(3775), vec(3773), vec(3772), vec(3770), vec(3768), vec(3767), vec(3765),
        vec(3763), vec(3761), vec(3760), vec(3758), vec(3756), vec(3755), vec(3753), vec(3751),
        vec(3749), vec(3748), vec(3746), vec(3744), vec(3742), vec(3741), vec(3739), vec(3737),
        vec(3735), vec(3733), vec(3732), vec(3730), vec(3728), vec(3726), vec(3724), vec(3723),
        vec(3721), vec(3719), vec(3717), vec(3715), vec(3714), vec(3712), vec(3710), vec(3708),
        vec(3706), vec(3704), vec(3703), vec(3701), vec(3699), vec(3697), vec(3695), vec(3693),
        vec(3691), vec(3690), vec(3688), vec(3686), vec(3684), vec(3682), vec(3680), vec(3678),
        vec(3676), vec(3674), vec(3672), vec(3671), vec(3669), vec(3667), vec(3665), vec(3663),
        vec(3661), vec(3659), vec(3657), vec(3655), vec(3653), vec(3651), vec(3649), vec(3647),
        vec(3645), vec(3643), vec(3641), vec(3639), vec(3637), vec(3635), vec(3634), vec(3632),
        vec(3630), vec(3628), vec(3626), vec(3624), vec(3622), vec(3620), vec(3617), vec(3615),
        vec(3613), vec(3611), vec(3609), vec(3607), vec(3605), vec(3603), vec(3601), vec(3599),
        vec(3597), vec(3595), vec(3593), vec(3591), vec(3589), vec(3587), vec(3585), vec(3583),
        vec(3581), vec(3579), vec(3576), vec(3574), vec(3572), vec(3570), vec(3568), vec(3566),
        vec(3564), vec(3562), vec(3560), vec(3557), vec(3555), vec(3553), vec(3551), vec(3549),
        vec(3547), vec(3545), vec(3543), vec(3540), vec(3538), vec(3536), vec(3534), vec(3532),
        vec(3530), vec(3527), vec(3525), vec(3523), vec(3521), vec(3519), vec(3517), vec(3514),
        vec(3512), vec(3510), vec(3508), vec(3506), vec(3503), vec(3501), vec(3499), vec(3497),
        vec(3494), vec(3492), vec(3490), vec(3488), vec(3486), vec(3483), vec(3481), vec(3479),
        vec(3477), vec(3474), vec(3472), vec(3470), vec(3468), vec(3465), vec(3463), vec(3461),
        vec(3458), vec(3456), vec(3454), vec(3452), vec(3449), vec(3447), vec(3445), vec(3442),
        vec(3440), vec(3438), vec(3436), vec(3433), vec(3431), vec(3429), vec(3426), vec(3424),
        vec(3422), vec(3419), vec(3417), vec(3415), vec(3412), vec(3410), vec(3408), vec(3405),
        vec(3403), vec(3401), vec(3398), vec(3396), vec(3393), vec(3391), vec(3389), vec(3386),
        vec(3384), vec(3382), vec(3379), vec(3377), vec(3374), vec(3372), vec(3370), vec(3367),
        vec(3365), vec(3362), vec(3360), vec(3358), vec(3355), vec(3353), vec(3350), vec(3348),
        vec(3345), vec(3343), vec(3341), vec(3338), vec(3336), vec(3333), vec(3331), vec(3328),
        vec(3326), vec(3323), vec(3321), vec(3319), vec(3316), vec(3314), vec(3311), vec(3309),
        vec(3306), vec(3304), vec(3301), vec(3299), vec(3296), vec(3294), vec(3291), vec(3289),
        vec(3286), vec(3284), vec(3281), vec(3279), vec(3276), vec(3274), vec(3271), vec(3269),
        vec(3266), vec(3264), vec(3261), vec(3259), vec(3256), vec(3254), vec(3251), vec(3248),
        vec(3246), vec(3243), vec(3241), vec(3238), vec(3236), vec(3233), vec(3231), vec(3228),
        vec(3225), vec(3223), vec(3220), vec(3218), vec(3215), vec(3213), vec(3210), vec(3207),
        vec(3205), vec(3202), vec(3200), vec(3197), vec(3194), vec(3192), vec(3189), vec(3187),
        vec(3184), vec(3181), vec(3179), vec(3176), vec(3173), vec(3171), vec(3168), vec(3166),
        vec(3163), vec(3160), vec(3158), vec(3155), vec(3152), vec(3150), vec(3147), vec(3144),
        vec(3142), vec(3139), vec(3137), vec(3134), vec(3131), vec(3129), vec(3126), vec(3123),
        vec(3120), vec(3118), vec(3115), vec(3112), vec(3110), vec(3107), vec(3104), vec(3102),
        vec(3099), vec(3096), vec(3094), vec(3091), vec(3088), vec(3086), vec(3083), vec(3080),
        vec(3077), vec(3075), vec(3072), vec(3069), vec(3066), vec(3064), vec(3061), vec(3058),
        vec(3056), vec(3053), vec(3050), vec(3047), vec(3045), vec(3042), vec(3039), vec(3036),
        vec(3034), vec(3031), vec(3028), vec(3025), vec(3023), vec(3020), vec(3017), vec(3014),
        vec(3012), vec(3009), vec(3006), vec(3003), vec(3000), vec(2998), vec(2995), vec(2992),
        vec(2989), vec(2986), vec(2984), vec(2981), vec(2978), vec(2975), vec(2972), vec(2970),
        vec(2967), vec(2964), vec(2961), vec(2958), vec(2956), vec(2953), vec(2950), vec(2947),
        vec(2944), vec(2942), vec(2939), vec(2936), vec(2933), vec(2930), vec(2927), vec(2925),
        vec(2922), vec(2919), vec(2916), vec(2913), vec(2910), vec(2907), vec(2905), vec(2902),
        vec(2899), vec(2896), vec(2893), vec(2890), vec(2887), vec(2885), vec(2882), vec(2879),
        vec(2876), vec(2873), vec(2870), vec(2867), vec(2864), vec(2862), vec(2859), vec(2856),
        vec(2853), vec(2850), vec(2847), vec(2844), vec(2841), vec(2838), vec(2836), vec(2833),
        vec(2830), vec(2827), vec(2824), vec(2821), vec(2818), vec(2815), vec(2812), vec(2809),
        vec(2806), vec(2804), vec(2801), vec(2798), vec(2795), vec(2792), vec(2789), vec(2786),
        vec(2783), vec(2780), vec(2777), vec(2774), vec(2771), vec(2768), vec(2765), vec(2763),
        vec(2760), vec(2757), vec(2754), vec(2751), vec(2748), vec(2745), vec(2742), vec(2739),
        vec(2736), vec(2733), vec(2730), vec(2727), vec(2724), vec(2721), vec(2718), vec(2715),
        vec(2712), vec(2709), vec(2706), vec(2703), vec(2700), vec(2697), vec(2694), vec(2691),
        vec(2688), vec(2685), vec(2682), vec(2679), vec(2676), vec(2673), vec(2670), vec(2668),
        vec(2665), vec(2662), vec(2659), vec(2656), vec(2653), vec(2650), vec(2647), vec(2644),
        vec(2640), vec(2637), vec(2634), vec(2631), vec(2628), vec(2625), vec(2622), vec(2619),
        vec(2616), vec(2613), vec(2610), vec(2607), vec(2604), vec(2601), vec(2598), vec(2595),
        vec(2592), vec(2589), vec(2586), vec(2583), vec(2580), vec(2577), vec(2574), vec(2571),
        vec(2568), vec(2565), vec(2562), vec(2559), vec(2556), vec(2553), vec(2550), vec(2547),
        vec(2544), vec(2541), vec(2537), vec(2534), vec(2531), vec(2528), vec(2525), vec(2522),
        vec(2519), vec(2516), vec(2513), vec(2510), vec(2507), vec(2504), vec(2501), vec(2498),
        vec(2495), vec(2492), vec(2489), vec(2485), vec(2482), vec(2479), vec(2476), vec(2473),
        vec(2470), vec(2467), vec(2464), vec(2461), vec(2458), vec(2455), vec(2452), vec(2449),
        vec(2446), vec(2442), vec(2439), vec(2436), vec(2433), vec(2430), vec(2427), vec(2424),
        vec(2421), vec(2418), vec(2415), vec(2412), vec(2408), vec(2405), vec(2402), vec(2399),
        vec(2396), vec(2393), vec(2390), vec(2387), vec(2384), vec(2381), vec(2377), vec(2374),
        vec(2371), vec(2368), vec(2365), vec(2362), vec(2359), vec(2356), vec(2353), vec(2350),
        vec(2346), vec(2343), vec(2340), vec(2337), vec(2334), vec(2331), vec(2328), vec(2325),
        vec(2322), vec(2318), vec(2315), vec(2312), vec(2309), vec(2306), vec(2303), vec(2300),
        vec(2297), vec(2294), vec(2290), vec(2287), vec(2284), vec(2281), vec(2278), vec(2275),
        vec(2272), vec(2269), vec(2265), vec(2262), vec(2259), vec(2256), vec(2253), vec(2250),
        vec(2247), vec(2244), vec(2240), vec(2237), vec(2234), vec(2231), vec(2228), vec(2225),
        vec(2222), vec(2219), vec(2215), vec(2212), vec(2209), vec(2206), vec(2203), vec(2200),
        vec(2197), vec(2193), vec(2190), vec(2187), vec(2184), vec(2181), vec(2178), vec(2175),
        vec(2172), vec(2168), vec(2165), vec(2162), vec(2159), vec(2156), vec(2153), vec(2150),
        vec(2146), vec(2143), vec(2140), vec(2137), vec(2134), vec(2131), vec(2128), vec(2124),
        vec(2121), vec(2118), vec(2115), vec(2112), vec(2109), vec(2106), vec(2102), vec(2099),
        vec(2096), vec(2093), vec(2090), vec(2087), vec(2084), vec(2080), vec(2077), vec(2074),
        vec(2071), vec(2068), vec(2065), vec(2062), vec(2058), vec(2055), vec(2052), vec(2049),
        vec(2046), vec(2043), vec(2040), vec(2037), vec(2033), vec(2030), vec(2027), vec(2024),
        vec(2021), vec(2018), vec(2015), vec(2011), vec(2008), vec(2005), vec(2002), vec(1999),
        vec(1996), vec(1993), vec(1989), vec(1986), vec(1983), vec(1980), vec(1977), vec(1974),
        vec(1971), vec(1967), vec(1964), vec(1961), vec(1958), vec(1955), vec(1952), vec(1949),
        vec(1945), vec(1942), vec(1939), vec(1936), vec(1933), vec(1930), vec(1927), vec(1923),
        vec(1920), vec(1917), vec(1914), vec(1911), vec(1908), vec(1905), vec(1902), vec(1898),
        vec(1895), vec(1892), vec(1889), vec(1886), vec(1883), vec(1880), vec(1876), vec(1873),
        vec(1870), vec(1867), vec(1864), vec(1861), vec(1858), vec(1855), vec(1851), vec(1848),
        vec(1845), vec(1842), vec(1839), vec(1836), vec(1833), vec(1830), vec(1826), vec(1823),
        vec(1820), vec(1817), vec(1814), vec(1811), vec(1808), vec(1805), vec(1801), vec(1798),
        vec(1795), vec(1792), vec(1789), vec(1786), vec(1783), vec(1780), vec(1777), vec(1773),
        vec(1770), vec(1767), vec(1764), vec(1761), vec(1758), vec(1755), vec(1752), vec(1749),
        vec(1745), vec(1742), vec(1739), vec(1736), vec(1733), vec(1730), vec(1727), vec(1724),
        vec(1721), vec(1718), vec(1714), vec(1711), vec(1708), vec(1705), vec(1702), vec(1699),
        vec(1696), vec(1693), vec(1690), vec(1687), vec(1683), vec(1680), vec(1677), vec(1674),
        vec(1671), vec(1668), vec(1665), vec(1662), vec(1659), vec(1656), vec(1653), vec(1649),
        vec(1646), vec(1643), vec(1640), vec(1637), vec(1634), vec(1631), vec(1628), vec(1625),
        vec(1622), vec(1619), vec(1616), vec(1613), vec(1610), vec(1606), vec(1603), vec(1600),
        vec(1597), vec(1594), vec(1591), vec(1588), vec(1585), vec(1582), vec(1579), vec(1576),
        vec(1573), vec(1570), vec(1567), vec(1564), vec(1561), vec(1558), vec(1554), vec(1551),
        vec(1548), vec(1545), vec(1542), vec(1539), vec(1536), vec(1533), vec(1530), vec(1527),
        vec(1524), vec(1521), vec(1518), vec(1515), vec(1512), vec(1509), vec(1506), vec(1503),
        vec(1500), vec(1497), vec(1494), vec(1491), vec(1488), vec(1485), vec(1482), vec(1479),
        vec(1476), vec(1473), vec(1470), vec(1467), vec(1464), vec(1461), vec(1458), vec(1455),
        vec(1451), vec(1448), vec(1445), vec(1442), vec(1439), vec(1436), vec(1433), vec(1430),
        vec(1427), vec(1425), vec(1422), vec(1419), vec(1416), vec(1413), vec(1410), vec(1407),
        vec(1404), vec(1401), vec(1398), vec(1395), vec(1392), vec(1389), vec(1386), vec(1383),
        vec(1380), vec(1377), vec(1374), vec(1371), vec(1368), vec(1365), vec(1362), vec(1359),
        vec(1356), vec(1353), vec(1350), vec(1347), vec(1344), vec(1341), vec(1338), vec(1335),
        vec(1332), vec(1330), vec(1327), vec(1324), vec(1321), vec(1318), vec(1315), vec(1312),
        vec(1309), vec(1306), vec(1303), vec(1300), vec(1297), vec(1294), vec(1291), vec(1289),
        vec(1286), vec(1283), vec(1280), vec(1277), vec(1274), vec(1271), vec(1268), vec(1265),
        vec(1262), vec(1259), vec(1257), vec(1254), vec(1251), vec(1248), vec(1245), vec(1242),
        vec(1239), vec(1236), vec(1233), vec(1231), vec(1228), vec(1225), vec(1222), vec(1219),
        vec(1216), vec(1213), vec(1210), vec(1208), vec(1205), vec(1202), vec(1199), vec(1196),
        vec(1193), vec(1190), vec(1188), vec(1185), vec(1182), vec(1179), vec(1176), vec(1173),
        vec(1170), vec(1168), vec(1165), vec(1162), vec(1159), vec(1156), vec(1153), vec(1151),
        vec(1148), vec(1145), vec(1142), vec(1139), vec(1137), vec(1134), vec(1131), vec(1128),
        vec(1125), vec(1123), vec(1120), vec(1117), vec(1114), vec(1111), vec(1109), vec(1106),
        vec(1103), vec(1100), vec(1097), vec(1095), vec(1092), vec(1089), vec(1086), vec(1083),
        vec(1081), vec(1078), vec(1075), vec(1072), vec(1070), vec(1067), vec(1064), vec(1061),
        vec(1059), vec(1056), vec(1053), vec(1050), vec(1048), vec(1045), vec(1042), vec(1039),
        vec(1037), vec(1034), vec(1031), vec(1029), vec(1026), vec(1023), vec(1020), vec(1018),
        vec(1015), vec(1012), vec(1009), vec(1007), vec(1004), vec(1001), vec(999), vec(996),
        vec(993), vec(991), vec(988), vec(985), vec(983), vec(980), vec(977), vec(975),
        vec(972), vec(969), vec(966), vec(964), vec(961), vec(958), vec(956), vec(953),
        vec(951), vec(948), vec(945), vec(943), vec(940), vec(937), vec(935), vec(932),
        vec(929), vec(927), vec(924), vec(922), vec(919), vec(916), vec(914), vec(911),
        vec(908), vec(906), vec(903), vec(901), vec(898), vec(895), vec(893), vec(890),
        vec(888), vec(885), vec(882), vec(880), vec(877), vec(875), vec(872), vec(870),
        vec(867), vec(864), vec(862), vec(859), vec(857), vec(854), vec(852), vec(849),
        vec(847), vec(844), vec(841), vec(839), vec(836), vec(834), vec(831), vec(829),
        vec(826), vec(824), vec(821), vec(819), vec(816), vec(814), vec(811), vec(809),
        vec(806), vec(804), vec(801), vec(799), vec(796), vec(794), vec(791), vec(789),
        vec(786), vec(784), vec(781), vec(779), vec(776), vec(774), vec(772), vec(769),
        vec(767), vec(764), vec(762), vec(759), vec(757), vec(754), vec(752), vec(750),
        vec(747), vec(745), vec(742), vec(740), vec(737), vec(735), vec(733), vec(730),
        vec(728), vec(725), vec(723), vec(721), vec(718), vec(716), vec(713), vec(711),
        vec(709), vec(706), vec(704), vec(702), vec(699), vec(697), vec(694), vec(692),
        vec(690), vec(687), vec(685), vec(683), vec(680), vec(678), vec(676), vec(673),
        vec(671), vec(669), vec(666), vec(664), vec(662), vec(659), vec(657), vec(655),
        vec(653), vec(650), vec(648), vec(646), vec(643), vec(641), vec(639), vec(637),
        vec(634), vec(632), vec(630), vec(627), vec(625), vec(623), vec(621), vec(618),
        vec(616), vec(614), vec(612), vec(609), vec(607), vec(605), vec(603), vec(601),
        vec(598), vec(596), vec(594), vec(592), vec(589), vec(587), vec(585), vec(583),
        vec(581), vec(578), vec(576), vec(574), vec(572), vec(570), vec(568), vec(565),
        vec(563), vec(561), vec(559), vec(557), vec(555), vec(552), vec(550), vec(548),
        vec(546), vec(544), vec(542), vec(540), vec(538), vec(535), vec(533), vec(531),
        vec(529), vec(527), vec(525), vec(523), vec(521), vec(519), vec(516), vec(514),
        vec(512), vec(510), vec(508), vec(506), vec(504), vec(502), vec(500), vec(498),
        vec(496), vec(494), vec(492), vec(490), vec(488), vec(486), vec(484), vec(482),
        vec(480), vec(478), vec(475), vec(473), vec(471), vec(469), vec(467), vec(465),
        vec(463), vec(461), vec(460), vec(458), vec(456), vec(454), vec(452), vec(450),
        vec(448), vec(446), vec(444), vec(442), vec(440), vec(438), vec(436), vec(434),
        vec(432), vec(430), vec(428), vec(426), vec(424), vec(423), vec(421), vec(419),
        vec(417), vec(415), vec(413), vec(411), vec(409), vec(407), vec(405), vec(404),
        vec(402), vec(400), vec(398), vec(396), vec(394), vec(392), vec(391), vec(389),
        vec(387), vec(385), vec(383), vec(381), vec(380), vec(378), vec(376), vec(374),
        vec(372), vec(371), vec(369), vec(367), vec(365), vec(363), vec(362), vec(360),
        vec(358), vec(356), vec(354), vec(353), vec(351), vec(349), vec(347), vec(346),
        vec(344), vec(342), vec(340), vec(339), vec(337), vec(335), vec(334), vec(332),
        vec(330), vec(328), vec(327), vec(325), vec(323), vec(322), vec(320), vec(318),
        vec(317), vec(315), vec(313), vec(312), vec(310), vec(308), vec(307), vec(305),
        vec(303), vec(302), vec(300), vec(298), vec(297), vec(295), vec(293), vec(292),
        vec(290), vec(289), vec(287), vec(285), vec(284), vec(282), vec(281), vec(279),
        vec(277), vec(276), vec(274), vec(273), vec(271), vec(270), vec(268), vec(267),
        vec(265), vec(263), vec(262), vec(260), vec(259), vec(257), vec(256), vec(254),
        vec(253), vec(251), vec(250), vec(248), vec(247), vec(245), vec(244), vec(242),
        vec(241), vec(239), vec(238), vec(236), vec(235), vec(233), vec(232), vec(231),
        vec(229), vec(228), vec(226), vec(225), vec(223), vec(222), vec(220), vec(219),
        vec(218), vec(216), vec(215), vec(213), vec(212), vec(211), vec(209), vec(208),
        vec(207), vec(205), vec(204), vec(202), vec(201), vec(200), vec(198), vec(197),
        vec(196), vec(194), vec(193), vec(192), vec(190), vec(189), vec(188), vec(186),
        vec(185), vec(184), vec(182), vec(181), vec(180), vec(179), vec(177), vec(176),
        vec(175), vec(174), vec(172), vec(171), vec(170), vec(168), vec(167), vec(166),
        vec(165), vec(164), vec(162), vec(161), vec(160), vec(159), vec(157), vec(156),
        vec(155), vec(154), vec(153), vec(151), vec(150), vec(149), vec(148), vec(147),
        vec(146), vec(144), vec(143), vec(142), vec(141), vec(140), vec(139), vec(138),
        vec(136), vec(135), vec(134), vec(133), vec(132), vec(131), vec(130), vec(129),
        vec(128), vec(126), vec(125), vec(124), vec(123), vec(122), vec(121), vec(120),
        vec(119), vec(118), vec(117), vec(116), vec(115), vec(114), vec(113), vec(112),
        vec(111), vec(110), vec(109), vec(108), vec(107), vec(106), vec(105), vec(104),
        vec(103), vec(102), vec(101), vec(100), vec(99), vec(98), vec(97), vec(96),
        vec(95), vec(94), vec(93), vec(92), vec(91), vec(90), vec(89), vec(88),
        vec(88), vec(87), vec(86), vec(85), vec(84), vec(83), vec(82), vec(81),
        vec(80), vec(80), vec(79), vec(78), vec(77), vec(76), vec(75), vec(74),
        vec(74), vec(73), vec(72), vec(71), vec(70), vec(69), vec(69), vec(68),
        vec(67), vec(66), vec(65), vec(65), vec(64), vec(63), vec(62), vec(62),
        vec(61), vec(60), vec(59), vec(59), vec(58), vec(57), vec(56), vec(56),
        vec(55), vec(54), vec(53), vec(53), vec(52), vec(51), vec(51), vec(50),
        vec(49), vec(49), vec(48), vec(47), vec(47), vec(46), vec(45), vec(45),
        vec(44), vec(43), vec(43), vec(42), vec(41), vec(41), vec(40), vec(40),
        vec(39), vec(38), vec(38), vec(37), vec(37), vec(36), vec(35), vec(35),
        vec(34), vec(34), vec(33), vec(32), vec(32), vec(31), vec(31), vec(30),
        vec(30), vec(29), vec(29), vec(28), vec(28), vec(27), vec(27), vec(26),
        vec(26), vec(25), vec(25), vec(24), vec(24), vec(23), vec(23), vec(22),
        vec(22), vec(21), vec(21), vec(20), vec(20), vec(20), vec(19), vec(19),
        vec(18), vec(18), vec(17), vec(17), vec(17), vec(16), vec(16), vec(16),
        vec(15), vec(15), vec(14), vec(14), vec(14), vec(13), vec(13), vec(13),
        vec(12), vec(12), vec(12), vec(11), vec(11), vec(11), vec(10), vec(10),
        vec(10), vec(9), vec(9), vec(9), vec(8), vec(8), vec(8), vec(8),
        vec(7), vec(7), vec(7), vec(7), vec(6), vec(6), vec(6), vec(6),
        vec(5), vec(5), vec(5), vec(5), vec(5), vec(4), vec(4), vec(4),
        vec(4), vec(4), vec(3), vec(3), vec(3), vec(3), vec(3), vec(3),
        vec(2), vec(2), vec(2), vec(2), vec(2), vec(2), vec(2), vec(1),
        vec(1), vec(1), vec(1), vec(1), vec(1), vec(1), vec(1), vec(1),
        vec(1), vec(0), vec(0), vec(0), vec(0), vec(0), vec(0), vec(0),
        vec(0), vec(0), vec(0), vec(0), vec(0), vec(0), vec(0), vec(0),
        vec(0), vec(0), vec(0), vec(0), vec(0), vec(0), vec(0), vec(0),
        vec(0), vec(0), vec(0), vec(0), vec(0), vec(0), vec(1), vec(1),
        vec(1), vec(1), vec(1), vec(1), vec(1), vec(1), vec(1), vec(1),
        vec(1), vec(2), vec(2), vec(2), vec(2), vec(2), vec(2), vec(2),
        vec(3), vec(3), vec(3), vec(3), vec(3), vec(3), vec(4), vec(4),
        vec(4), vec(4), vec(4), vec(5), vec(5), vec(5), vec(5), vec(5),
        vec(6), vec(6), vec(6), vec(6), vec(7), vec(7), vec(7), vec(7),
        vec(8), vec(8), vec(8), vec(9), vec(9), vec(9), vec(9), vec(10),
        vec(10), vec(10), vec(11), vec(11), vec(11), vec(12), vec(12), vec(12),
        vec(13), vec(13), vec(13), vec(14), vec(14), vec(15), vec(15), vec(15),
        vec(16), vec(16), vec(16), vec(17), vec(17), vec(18), vec(18), vec(19),
        vec(19), vec(19), vec(20), vec(20), vec(21), vec(21), vec(22), vec(22),
        vec(23), vec(23), vec(23), vec(24), vec(24), vec(25), vec(25), vec(26),
        vec(26), vec(27), vec(27), vec(28), vec(28), vec(29), vec(29), vec(30),
        vec(31), vec(31), vec(32), vec(32), vec(33), vec(33), vec(34), vec(34),
        vec(35), vec(36), vec(36), vec(37), vec(37), vec(38), vec(39), vec(39),
        vec(40), vec(40), vec(41), vec(42), vec(42), vec(43), vec(44), vec(44),
        vec(45), vec(46), vec(46), vec(47), vec(48), vec(48), vec(49), vec(50),
        vec(50), vec(51), vec(52), vec(52), vec(53), vec(54), vec(55), vec(55),
        vec(56), vec(57), vec(57), vec(58), vec(59), vec(60), vec(60), vec(61),
        vec(62), vec(63), vec(64), vec(64), vec(65), vec(66), vec(67), vec(67),
        vec(68), vec(69), vec(70), vec(71), vec(72), vec(72), vec(73), vec(74),
        vec(75), vec(76), vec(77), vec(77), vec(78), vec(79), vec(80), vec(81),
        vec(82), vec(83), vec(83), vec(84), vec(85), vec(86), vec(87), vec(88),
        vec(89), vec(90), vec(91), vec(92), vec(93), vec(94), vec(94), vec(95),
        vec(96), vec(97), vec(98), vec(99), vec(100), vec(101), vec(102), vec(103),
        vec(104), vec(105), vec(106), vec(107), vec(108), vec(109), vec(110), vec(111),
        vec(112), vec(113), vec(114), vec(115), vec(116), vec(117), vec(118), vec(119),
        vec(121), vec(122), vec(123), vec(124), vec(125), vec(126), vec(127), vec(128),
        vec(129), vec(130), vec(131), vec(132), vec(134), vec(135), vec(136), vec(137),
        vec(138), vec(139), vec(140), vec(142), vec(143), vec(144), vec(145), vec(146),
        vec(147), vec(149), vec(150), vec(151), vec(152), vec(153), vec(154), vec(156),
        vec(157), vec(158), vec(159), vec(160), vec(162), vec(163), vec(164), vec(165),
        vec(167), vec(168), vec(169), vec(170), vec(172), vec(173), vec(174), vec(175),
        vec(177), vec(178), vec(179), vec(181), vec(182), vec(183), vec(184), vec(186),
        vec(187), vec(188), vec(190), vec(191), vec(192), vec(194), vec(195), vec(196),
        vec(198), vec(199), vec(200), vec(202), vec(203), vec(204), vec(206), vec(207),
        vec(209), vec(210), vec(211), vec(213), vec(214), vec(216), vec(217), vec(218),
        vec(220), vec(221), vec(223), vec(224), vec(225), vec(227), vec(228), vec(230),
        vec(231), vec(233), vec(234), vec(236), vec(237), vec(239), vec(240), vec(242),
        vec(243), vec(244), vec(246), vec(247), vec(249), vec(250), vec(252), vec(253),
        vec(255), vec(257), vec(258), vec(260), vec(261), vec(263), vec(264), vec(266),
        vec(267), vec(269), vec(270), vec(272), vec(274), vec(275), vec(277), vec(278),
        vec(280), vec(281), vec(283), vec(285), vec(286), vec(288), vec(289), vec(291),
        vec(293), vec(294), vec(296), vec(298), vec(299), vec(301), vec(302), vec(304),
        vec(306), vec(307), vec(309), vec(311), vec(312), vec(314), vec(316), vec(317),
        vec(319), vec(321), vec(322), vec(324), vec(326), vec(328), vec(329), vec(331),
        vec(333), vec(334), vec(336), vec(338), vec(340), vec(341), vec(343), vec(345),
        vec(347), vec(348), vec(350), vec(352), vec(354), vec(355), vec(357), vec(359),
        vec(361), vec(362), vec(364), vec(366), vec(368), vec(370), vec(371), vec(373),
        vec(375), vec(377), vec(379), vec(380), vec(382), vec(384), vec(386), vec(388),
        vec(390), vec(391), vec(393), vec(395), vec(397), vec(399), vec(401), vec(403),
        vec(405), vec(406), vec(408), vec(410), vec(412), vec(414), vec(416), vec(418),
        vec(420), vec(422), vec(423), vec(425), vec(427), vec(429), vec(431), vec(433),
        vec(435), vec(437), vec(439), vec(441), vec(443), vec(445), vec(447), vec(449),
        vec(451), vec(453), vec(455), vec(457), vec(459), vec(461), vec(462), vec(464),
        vec(466), vec(468), vec(470), vec(472), vec(474), vec(477), vec(479), vec(481),
        vec(483), vec(485), vec(487), vec(489), vec(491), vec(493), vec(495), vec(497),
        vec(499), vec(501), vec(503), vec(505), vec(507), vec(509), vec(511), vec(513),
        vec(515), vec(518), vec(520), vec(522), vec(524), vec(526), vec(528), vec(530),
        vec(532), vec(534), vec(536), vec(539), vec(541), vec(543), vec(545), vec(547),
        vec(549), vec(551), vec(554), vec(556), vec(558), vec(560), vec(562), vec(564),
        vec(566), vec(569), vec(571), vec(573), vec(575), vec(577), vec(580), vec(582),
        vec(584), vec(586), vec(588), vec(591), vec(593), vec(595), vec(597), vec(599),
        vec(602), vec(604), vec(606), vec(608), vec(611), vec(613), vec(615), vec(617),
        vec(620), vec(622), vec(624), vec(626), vec(629), vec(631), vec(633), vec(635),
        vec(638), vec(640), vec(642), vec(645), vec(647), vec(649), vec(651), vec(654),
        vec(656), vec(658), vec(661), vec(663), vec(665), vec(668), vec(670), vec(672),
        vec(675), vec(677), vec(679), vec(682), vec(684), vec(686), vec(689), vec(691),
        vec(693), vec(696), vec(698), vec(700), vec(703), vec(705), vec(707), vec(710),
        vec(712), vec(715), vec(717), vec(719), vec(722), vec(724), vec(727), vec(729),
        vec(731), vec(734), vec(736), vec(739), vec(741), vec(743), vec(746), vec(748),
        vec(751), vec(753), vec(756), vec(758), vec(760), vec(763), vec(765), vec(768),
        vec(770), vec(773), vec(775), vec(778), vec(780), vec(783), vec(785), vec(788),
        vec(790), vec(793), vec(795), vec(797), vec(800), vec(802), vec(805), vec(807),
        vec(810), vec(812), vec(815), vec(817), vec(820), vec(823), vec(825), vec(828),
        vec(830), vec(833), vec(835), vec(838), vec(840), vec(843), vec(845), vec(848),
        vec(850), vec(853), vec(855), vec(858), vec(861), vec(863), vec(866), vec(868),
        vec(871), vec(873), vec(876), vec(879), vec(881), vec(884), vec(886), vec(889),
        vec(892), vec(894), vec(897), vec(899), vec(902), vec(905), vec(907), vec(910),
        vec(912), vec(915), vec(918), vec(920), vec(923), vec(925), vec(928), vec(931),
        vec(933), vec(936), vec(939), vec(941), vec(944), vec(947), vec(949), vec(952),
        vec(955), vec(957), vec(960), vec(962), vec(965), vec(968), vec(970), vec(973),
        vec(976), vec(979), vec(981), vec(984), vec(987), vec(989), vec(992), vec(995),
        vec(997), vec(1000), vec(1003), vec(1005), vec(1008), vec(1011), vec(1014), vec(1016),
        vec(1019), vec(1022), vec(1024), vec(1027), vec(1030), vec(1033), vec(1035), vec(1038),
        vec(1041), vec(1044), vec(1046), vec(1049), vec(1052), vec(1055), vec(1057), vec(1060),
        vec(1063), vec(1066), vec(1068), vec(1071), vec(1074), vec(1077), vec(1079), vec(1082),
        vec(1085), vec(1088), vec(1090), vec(1093), vec(1096), vec(1099), vec(1102), vec(1104),
        vec(1107), vec(1110), vec(1113), vec(1116), vec(1118), vec(1121), vec(1124), vec(1127),
        vec(1130), vec(1132), vec(1135), vec(1138), vec(1141), vec(1144), vec(1146), vec(1149),
        vec(1152), vec(1155), vec(1158), vec(1161), vec(1163), vec(1166), vec(1169), vec(1172),
        vec(1175), vec(1178), vec(1180), vec(1183), vec(1186), vec(1189), vec(1192), vec(1195),
        vec(1198), vec(1200), vec(1203), vec(1206), vec(1209), vec(1212), vec(1215), vec(1218),
        vec(1220), vec(1223), vec(1226), vec(1229), vec(1232), vec(1235), vec(1238), vec(1241),
        vec(1244), vec(1246), vec(1249), vec(1252), vec(1255), vec(1258), vec(1261), vec(1264),
        vec(1267), vec(1270), vec(1272), vec(1275), vec(1278), vec(1281), vec(1284), vec(1287),
        vec(1290), vec(1293), vec(1296), vec(1299), vec(1302), vec(1305), vec(1308), vec(1310),
        vec(1313), vec(1316), vec(1319), vec(1322), vec(1325), vec(1328), vec(1331), vec(1334),
        vec(1337), vec(1340), vec(1343), vec(1346), vec(1349), vec(1352), vec(1355), vec(1358),
        vec(1361), vec(1363), vec(1366), vec(1369), vec(1372), vec(1375), vec(1378), vec(1381),
        vec(1384), vec(1387), vec(1390), vec(1393), vec(1396), vec(1399), vec(1402), vec(1405),
        vec(1408), vec(1411), vec(1414), vec(1417), vec(1420), vec(1423), vec(1426), vec(1429),
        vec(1432), vec(1435), vec(1438), vec(1441), vec(1444), vec(1447), vec(1450), vec(1453),
        vec(1456), vec(1459), vec(1462), vec(1465), vec(1468), vec(1471), vec(1474), vec(1477),
        vec(1480), vec(1483), vec(1486), vec(1489), vec(1492), vec(1495), vec(1498), vec(1501),
        vec(1504), vec(1507), vec(1510), vec(1513), vec(1516), vec(1519), vec(1523), vec(1526),
        vec(1529), vec(1532), vec(1535), vec(1538), vec(1541), vec(1544), vec(1547), vec(1550),
        vec(1553), vec(1556), vec(1559), vec(1562), vec(1565), vec(1568), vec(1571), vec(1574),
        vec(1577), vec(1580), vec(1583), vec(1587), vec(1590), vec(1593), vec(1596), vec(1599),
        vec(1602), vec(1605), vec(1608), vec(1611), vec(1614), vec(1617), vec(1620), vec(1623),
        vec(1626), vec(1629), vec(1633), vec(1636), vec(1639), vec(1642), vec(1645), vec(1648),
        vec(1651), vec(1654), vec(1657), vec(1660), vec(1663), vec(1666), vec(1670), vec(1673),
        vec(1676), vec(1679), vec(1682), vec(1685), vec(1688), vec(1691), vec(1694), vec(1697),
        vec(1700), vec(1704), vec(1707), vec(1710), vec(1713), vec(1716), vec(1719), vec(1722),
        vec(1725), vec(1728), vec(1731), vec(1735), vec(1738), vec(1741), vec(1744), vec(1747),
        vec(1750), vec(1753), vec(1756), vec(1759), vec(1763), vec(1766), vec(1769), vec(1772),
        vec(1775), vec(1778), vec(1781), vec(1784), vec(1787), vec(1791), vec(1794), vec(1797),
        vec(1800), vec(1803), vec(1806), vec(1809), vec(1812), vec(1816), vec(1819), vec(1822),
        vec(1825), vec(1828), vec(1831), vec(1834), vec(1837), vec(1841), vec(1844), vec(1847),
        vec(1850), vec(1853), vec(1856), vec(1859), vec(1862), vec(1866), vec(1869), vec(1872),
        vec(1875), vec(1878), vec(1881), vec(1884), vec(1887), vec(1891), vec(1894), vec(1897),
        vec(1900), vec(1903), vec(1906), vec(1909), vec(1913), vec(1916), vec(1919), vec(1922),
        vec(1925), vec(1928), vec(1931), vec(1934), vec(1938), vec(1941), vec(1944), vec(1947),
        vec(1950), vec(1953), vec(1956), vec(1960), vec(1963), vec(1966), vec(1969), vec(1972),
        vec(1975), vec(1978), vec(1982), vec(1985), vec(1988), vec(1991), vec(1994), vec(1997),
        vec(2000), vec(2004), vec(2007), vec(2010), vec(2013), vec(2016), vec(2019), vec(2022),
        vec(2026), vec(2029), vec(2032), vec(2035), vec(2038), vec(2041), vec(2044), vec(2047)
    );

end package sin_1T_4096s_12b_pkg;

package body sin_1T_4096s_12b_pkg is

    function vec(value : integer) return std_logic_vector is
    begin
        return std_logic_vector(to_unsigned(value, 12));
    end function vec;

end package body sin_1T_4096s_12b_pkg;
