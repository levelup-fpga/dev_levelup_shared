-- Generated curve samples
-- ==================================================
-- Y_real values (no virtual zoom)
-- Curve type: sin
-- Number of samples: 2048
-- Bit range: 12 bits (0 to 4095)
-- ==================================================

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

package sin_1T_2048s_12b_pkg is

    type sample_array_t is array (0 to 2047) of std_logic_vector(11 downto 0);

    function vec(value : integer) return std_logic_vector;

    constant SAMPLES : sample_array_t := (
        vec(2048), vec(2054), vec(2060), vec(2066), vec(2073), vec(2079), vec(2085), vec(2091),
        vec(2098), vec(2104), vec(2110), vec(2117), vec(2123), vec(2129), vec(2135), vec(2142),
        vec(2148), vec(2154), vec(2161), vec(2167), vec(2173), vec(2179), vec(2186), vec(2192),
        vec(2198), vec(2204), vec(2211), vec(2217), vec(2223), vec(2230), vec(2236), vec(2242),
        vec(2248), vec(2255), vec(2261), vec(2267), vec(2273), vec(2280), vec(2286), vec(2292),
        vec(2298), vec(2304), vec(2311), vec(2317), vec(2323), vec(2329), vec(2336), vec(2342),
        vec(2348), vec(2354), vec(2361), vec(2367), vec(2373), vec(2379), vec(2385), vec(2392),
        vec(2398), vec(2404), vec(2410), vec(2416), vec(2422), vec(2429), vec(2435), vec(2441),
        vec(2447), vec(2453), vec(2459), vec(2466), vec(2472), vec(2478), vec(2484), vec(2490),
        vec(2496), vec(2502), vec(2509), vec(2515), vec(2521), vec(2527), vec(2533), vec(2539),
        vec(2545), vec(2551), vec(2557), vec(2564), vec(2570), vec(2576), vec(2582), vec(2588),
        vec(2594), vec(2600), vec(2606), vec(2612), vec(2618), vec(2624), vec(2630), vec(2636),
        vec(2642), vec(2648), vec(2654), vec(2660), vec(2666), vec(2672), vec(2678), vec(2684),
        vec(2690), vec(2696), vec(2702), vec(2708), vec(2714), vec(2720), vec(2726), vec(2732),
        vec(2738), vec(2744), vec(2749), vec(2755), vec(2761), vec(2767), vec(2773), vec(2779),
        vec(2785), vec(2791), vec(2796), vec(2802), vec(2808), vec(2814), vec(2820), vec(2826),
        vec(2831), vec(2837), vec(2843), vec(2849), vec(2855), vec(2860), vec(2866), vec(2872),
        vec(2878), vec(2883), vec(2889), vec(2895), vec(2901), vec(2906), vec(2912), vec(2918),
        vec(2923), vec(2929), vec(2935), vec(2940), vec(2946), vec(2952), vec(2957), vec(2963),
        vec(2968), vec(2974), vec(2980), vec(2985), vec(2991), vec(2996), vec(3002), vec(3008),
        vec(3013), vec(3019), vec(3024), vec(3030), vec(3035), vec(3041), vec(3046), vec(3052),
        vec(3057), vec(3063), vec(3068), vec(3074), vec(3079), vec(3084), vec(3090), vec(3095),
        vec(3101), vec(3106), vec(3111), vec(3117), vec(3122), vec(3127), vec(3133), vec(3138),
        vec(3143), vec(3149), vec(3154), vec(3159), vec(3165), vec(3170), vec(3175), vec(3180),
        vec(3186), vec(3191), vec(3196), vec(3201), vec(3206), vec(3212), vec(3217), vec(3222),
        vec(3227), vec(3232), vec(3237), vec(3242), vec(3247), vec(3253), vec(3258), vec(3263),
        vec(3268), vec(3273), vec(3278), vec(3283), vec(3288), vec(3293), vec(3298), vec(3303),
        vec(3308), vec(3313), vec(3318), vec(3323), vec(3327), vec(3332), vec(3337), vec(3342),
        vec(3347), vec(3352), vec(3357), vec(3361), vec(3366), vec(3371), vec(3376), vec(3381),
        vec(3385), vec(3390), vec(3395), vec(3400), vec(3404), vec(3409), vec(3414), vec(3418),
        vec(3423), vec(3428), vec(3432), vec(3437), vec(3442), vec(3446), vec(3451), vec(3455),
        vec(3460), vec(3464), vec(3469), vec(3473), vec(3478), vec(3482), vec(3487), vec(3491),
        vec(3496), vec(3500), vec(3505), vec(3509), vec(3514), vec(3518), vec(3522), vec(3527),
        vec(3531), vec(3535), vec(3540), vec(3544), vec(3548), vec(3552), vec(3557), vec(3561),
        vec(3565), vec(3569), vec(3574), vec(3578), vec(3582), vec(3586), vec(3590), vec(3594),
        vec(3598), vec(3603), vec(3607), vec(3611), vec(3615), vec(3619), vec(3623), vec(3627),
        vec(3631), vec(3635), vec(3639), vec(3643), vec(3647), vec(3651), vec(3654), vec(3658),
        vec(3662), vec(3666), vec(3670), vec(3674), vec(3678), vec(3681), vec(3685), vec(3689),
        vec(3693), vec(3696), vec(3700), vec(3704), vec(3707), vec(3711), vec(3715), vec(3718),
        vec(3722), vec(3726), vec(3729), vec(3733), vec(3736), vec(3740), vec(3743), vec(3747),
        vec(3750), vec(3754), vec(3757), vec(3761), vec(3764), vec(3768), vec(3771), vec(3775),
        vec(3778), vec(3781), vec(3785), vec(3788), vec(3791), vec(3794), vec(3798), vec(3801),
        vec(3804), vec(3807), vec(3811), vec(3814), vec(3817), vec(3820), vec(3823), vec(3826),
        vec(3830), vec(3833), vec(3836), vec(3839), vec(3842), vec(3845), vec(3848), vec(3851),
        vec(3854), vec(3857), vec(3860), vec(3863), vec(3865), vec(3868), vec(3871), vec(3874),
        vec(3877), vec(3880), vec(3882), vec(3885), vec(3888), vec(3891), vec(3893), vec(3896),
        vec(3899), vec(3902), vec(3904), vec(3907), vec(3909), vec(3912), vec(3915), vec(3917),
        vec(3920), vec(3922), vec(3925), vec(3927), vec(3930), vec(3932), vec(3935), vec(3937),
        vec(3940), vec(3942), vec(3944), vec(3947), vec(3949), vec(3951), vec(3954), vec(3956),
        vec(3958), vec(3960), vec(3963), vec(3965), vec(3967), vec(3969), vec(3971), vec(3974),
        vec(3976), vec(3978), vec(3980), vec(3982), vec(3984), vec(3986), vec(3988), vec(3990),
        vec(3992), vec(3994), vec(3996), vec(3998), vec(4000), vec(4002), vec(4004), vec(4005),
        vec(4007), vec(4009), vec(4011), vec(4013), vec(4014), vec(4016), vec(4018), vec(4019),
        vec(4021), vec(4023), vec(4024), vec(4026), vec(4028), vec(4029), vec(4031), vec(4032),
        vec(4034), vec(4035), vec(4037), vec(4038), vec(4040), vec(4041), vec(4043), vec(4044),
        vec(4046), vec(4047), vec(4048), vec(4050), vec(4051), vec(4052), vec(4053), vec(4055),
        vec(4056), vec(4057), vec(4058), vec(4060), vec(4061), vec(4062), vec(4063), vec(4064),
        vec(4065), vec(4066), vec(4067), vec(4068), vec(4069), vec(4070), vec(4071), vec(4072),
        vec(4073), vec(4074), vec(4075), vec(4076), vec(4077), vec(4077), vec(4078), vec(4079),
        vec(4080), vec(4081), vec(4081), vec(4082), vec(4083), vec(4083), vec(4084), vec(4085),
        vec(4085), vec(4086), vec(4086), vec(4087), vec(4088), vec(4088), vec(4089), vec(4089),
        vec(4090), vec(4090), vec(4090), vec(4091), vec(4091), vec(4092), vec(4092), vec(4092),
        vec(4093), vec(4093), vec(4093), vec(4093), vec(4094), vec(4094), vec(4094), vec(4094),
        vec(4094), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095),
        vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4095), vec(4094),
        vec(4094), vec(4094), vec(4094), vec(4094), vec(4094), vec(4093), vec(4093), vec(4093),
        vec(4092), vec(4092), vec(4092), vec(4091), vec(4091), vec(4091), vec(4090), vec(4090),
        vec(4089), vec(4089), vec(4088), vec(4088), vec(4087), vec(4087), vec(4086), vec(4086),
        vec(4085), vec(4084), vec(4084), vec(4083), vec(4082), vec(4082), vec(4081), vec(4080),
        vec(4079), vec(4079), vec(4078), vec(4077), vec(4076), vec(4075), vec(4074), vec(4074),
        vec(4073), vec(4072), vec(4071), vec(4070), vec(4069), vec(4068), vec(4067), vec(4066),
        vec(4065), vec(4063), vec(4062), vec(4061), vec(4060), vec(4059), vec(4058), vec(4057),
        vec(4055), vec(4054), vec(4053), vec(4052), vec(4050), vec(4049), vec(4048), vec(4046),
        vec(4045), vec(4043), vec(4042), vec(4041), vec(4039), vec(4038), vec(4036), vec(4035),
        vec(4033), vec(4032), vec(4030), vec(4029), vec(4027), vec(4025), vec(4024), vec(4022),
        vec(4020), vec(4019), vec(4017), vec(4015), vec(4013), vec(4012), vec(4010), vec(4008),
        vec(4006), vec(4004), vec(4003), vec(4001), vec(3999), vec(3997), vec(3995), vec(3993),
        vec(3991), vec(3989), vec(3987), vec(3985), vec(3983), vec(3981), vec(3979), vec(3977),
        vec(3975), vec(3973), vec(3970), vec(3968), vec(3966), vec(3964), vec(3962), vec(3959),
        vec(3957), vec(3955), vec(3953), vec(3950), vec(3948), vec(3946), vec(3943), vec(3941),
        vec(3938), vec(3936), vec(3934), vec(3931), vec(3929), vec(3926), vec(3924), vec(3921),
        vec(3919), vec(3916), vec(3913), vec(3911), vec(3908), vec(3906), vec(3903), vec(3900),
        vec(3898), vec(3895), vec(3892), vec(3889), vec(3887), vec(3884), vec(3881), vec(3878),
        vec(3875), vec(3873), vec(3870), vec(3867), vec(3864), vec(3861), vec(3858), vec(3855),
        vec(3852), vec(3849), vec(3846), vec(3843), vec(3840), vec(3837), vec(3834), vec(3831),
        vec(3828), vec(3825), vec(3822), vec(3819), vec(3815), vec(3812), vec(3809), vec(3806),
        vec(3803), vec(3799), vec(3796), vec(3793), vec(3790), vec(3786), vec(3783), vec(3780),
        vec(3776), vec(3773), vec(3769), vec(3766), vec(3763), vec(3759), vec(3756), vec(3752),
        vec(3749), vec(3745), vec(3742), vec(3738), vec(3735), vec(3731), vec(3727), vec(3724),
        vec(3720), vec(3717), vec(3713), vec(3709), vec(3706), vec(3702), vec(3698), vec(3694),
        vec(3691), vec(3687), vec(3683), vec(3679), vec(3676), vec(3672), vec(3668), vec(3664),
        vec(3660), vec(3656), vec(3652), vec(3649), vec(3645), vec(3641), vec(3637), vec(3633),
        vec(3629), vec(3625), vec(3621), vec(3617), vec(3613), vec(3609), vec(3605), vec(3600),
        vec(3596), vec(3592), vec(3588), vec(3584), vec(3580), vec(3576), vec(3571), vec(3567),
        vec(3563), vec(3559), vec(3555), vec(3550), vec(3546), vec(3542), vec(3537), vec(3533),
        vec(3529), vec(3524), vec(3520), vec(3516), vec(3511), vec(3507), vec(3503), vec(3498),
        vec(3494), vec(3489), vec(3485), vec(3480), vec(3476), vec(3471), vec(3467), vec(3462),
        vec(3458), vec(3453), vec(3448), vec(3444), vec(3439), vec(3435), vec(3430), vec(3425),
        vec(3421), vec(3416), vec(3411), vec(3407), vec(3402), vec(3397), vec(3393), vec(3388),
        vec(3383), vec(3378), vec(3373), vec(3369), vec(3364), vec(3359), vec(3354), vec(3349),
        vec(3345), vec(3340), vec(3335), vec(3330), vec(3325), vec(3320), vec(3315), vec(3310),
        vec(3305), vec(3300), vec(3295), vec(3290), vec(3285), vec(3280), vec(3275), vec(3270),
        vec(3265), vec(3260), vec(3255), vec(3250), vec(3245), vec(3240), vec(3235), vec(3230),
        vec(3224), vec(3219), vec(3214), vec(3209), vec(3204), vec(3199), vec(3193), vec(3188),
        vec(3183), vec(3178), vec(3172), vec(3167), vec(3162), vec(3157), vec(3151), vec(3146),
        vec(3141), vec(3135), vec(3130), vec(3125), vec(3119), vec(3114), vec(3109), vec(3103),
        vec(3098), vec(3092), vec(3087), vec(3082), vec(3076), vec(3071), vec(3065), vec(3060),
        vec(3054), vec(3049), vec(3043), vec(3038), vec(3032), vec(3027), vec(3021), vec(3016),
        vec(3010), vec(3005), vec(2999), vec(2994), vec(2988), vec(2983), vec(2977), vec(2971),
        vec(2966), vec(2960), vec(2954), vec(2949), vec(2943), vec(2937), vec(2932), vec(2926),
        vec(2920), vec(2915), vec(2909), vec(2903), vec(2898), vec(2892), vec(2886), vec(2880),
        vec(2875), vec(2869), vec(2863), vec(2857), vec(2852), vec(2846), vec(2840), vec(2834),
        vec(2829), vec(2823), vec(2817), vec(2811), vec(2805), vec(2799), vec(2794), vec(2788),
        vec(2782), vec(2776), vec(2770), vec(2764), vec(2758), vec(2752), vec(2746), vec(2741),
        vec(2735), vec(2729), vec(2723), vec(2717), vec(2711), vec(2705), vec(2699), vec(2693),
        vec(2687), vec(2681), vec(2675), vec(2669), vec(2663), vec(2657), vec(2651), vec(2645),
        vec(2639), vec(2633), vec(2627), vec(2621), vec(2615), vec(2609), vec(2603), vec(2597),
        vec(2591), vec(2585), vec(2579), vec(2573), vec(2567), vec(2560), vec(2554), vec(2548),
        vec(2542), vec(2536), vec(2530), vec(2524), vec(2518), vec(2512), vec(2506), vec(2499),
        vec(2493), vec(2487), vec(2481), vec(2475), vec(2469), vec(2463), vec(2456), vec(2450),
        vec(2444), vec(2438), vec(2432), vec(2426), vec(2419), vec(2413), vec(2407), vec(2401),
        vec(2395), vec(2388), vec(2382), vec(2376), vec(2370), vec(2364), vec(2357), vec(2351),
        vec(2345), vec(2339), vec(2333), vec(2326), vec(2320), vec(2314), vec(2308), vec(2301),
        vec(2295), vec(2289), vec(2283), vec(2276), vec(2270), vec(2264), vec(2258), vec(2251),
        vec(2245), vec(2239), vec(2233), vec(2226), vec(2220), vec(2214), vec(2208), vec(2201),
        vec(2195), vec(2189), vec(2183), vec(2176), vec(2170), vec(2164), vec(2157), vec(2151),
        vec(2145), vec(2139), vec(2132), vec(2126), vec(2120), vec(2113), vec(2107), vec(2101),
        vec(2095), vec(2088), vec(2082), vec(2076), vec(2069), vec(2063), vec(2057), vec(2051),
        vec(2044), vec(2038), vec(2032), vec(2026), vec(2019), vec(2013), vec(2007), vec(2000),
        vec(1994), vec(1988), vec(1982), vec(1975), vec(1969), vec(1963), vec(1956), vec(1950),
        vec(1944), vec(1938), vec(1931), vec(1925), vec(1919), vec(1912), vec(1906), vec(1900),
        vec(1894), vec(1887), vec(1881), vec(1875), vec(1869), vec(1862), vec(1856), vec(1850),
        vec(1844), vec(1837), vec(1831), vec(1825), vec(1819), vec(1812), vec(1806), vec(1800),
        vec(1794), vec(1787), vec(1781), vec(1775), vec(1769), vec(1762), vec(1756), vec(1750),
        vec(1744), vec(1738), vec(1731), vec(1725), vec(1719), vec(1713), vec(1707), vec(1700),
        vec(1694), vec(1688), vec(1682), vec(1676), vec(1669), vec(1663), vec(1657), vec(1651),
        vec(1645), vec(1639), vec(1632), vec(1626), vec(1620), vec(1614), vec(1608), vec(1602),
        vec(1596), vec(1589), vec(1583), vec(1577), vec(1571), vec(1565), vec(1559), vec(1553),
        vec(1547), vec(1541), vec(1535), vec(1528), vec(1522), vec(1516), vec(1510), vec(1504),
        vec(1498), vec(1492), vec(1486), vec(1480), vec(1474), vec(1468), vec(1462), vec(1456),
        vec(1450), vec(1444), vec(1438), vec(1432), vec(1426), vec(1420), vec(1414), vec(1408),
        vec(1402), vec(1396), vec(1390), vec(1384), vec(1378), vec(1372), vec(1366), vec(1360),
        vec(1354), vec(1349), vec(1343), vec(1337), vec(1331), vec(1325), vec(1319), vec(1313),
        vec(1307), vec(1301), vec(1296), vec(1290), vec(1284), vec(1278), vec(1272), vec(1266),
        vec(1261), vec(1255), vec(1249), vec(1243), vec(1238), vec(1232), vec(1226), vec(1220),
        vec(1215), vec(1209), vec(1203), vec(1197), vec(1192), vec(1186), vec(1180), vec(1175),
        vec(1169), vec(1163), vec(1158), vec(1152), vec(1146), vec(1141), vec(1135), vec(1129),
        vec(1124), vec(1118), vec(1112), vec(1107), vec(1101), vec(1096), vec(1090), vec(1085),
        vec(1079), vec(1074), vec(1068), vec(1063), vec(1057), vec(1052), vec(1046), vec(1041),
        vec(1035), vec(1030), vec(1024), vec(1019), vec(1013), vec(1008), vec(1003), vec(997),
        vec(992), vec(986), vec(981), vec(976), vec(970), vec(965), vec(960), vec(954),
        vec(949), vec(944), vec(938), vec(933), vec(928), vec(923), vec(917), vec(912),
        vec(907), vec(902), vec(896), vec(891), vec(886), vec(881), vec(876), vec(871),
        vec(865), vec(860), vec(855), vec(850), vec(845), vec(840), vec(835), vec(830),
        vec(825), vec(820), vec(815), vec(810), vec(805), vec(800), vec(795), vec(790),
        vec(785), vec(780), vec(775), vec(770), vec(765), vec(760), vec(755), vec(750),
        vec(746), vec(741), vec(736), vec(731), vec(726), vec(722), vec(717), vec(712),
        vec(707), vec(702), vec(698), vec(693), vec(688), vec(684), vec(679), vec(674),
        vec(670), vec(665), vec(660), vec(656), vec(651), vec(647), vec(642), vec(637),
        vec(633), vec(628), vec(624), vec(619), vec(615), vec(610), vec(606), vec(601),
        vec(597), vec(592), vec(588), vec(584), vec(579), vec(575), vec(571), vec(566),
        vec(562), vec(558), vec(553), vec(549), vec(545), vec(540), vec(536), vec(532),
        vec(528), vec(524), vec(519), vec(515), vec(511), vec(507), vec(503), vec(499),
        vec(495), vec(490), vec(486), vec(482), vec(478), vec(474), vec(470), vec(466),
        vec(462), vec(458), vec(454), vec(450), vec(446), vec(443), vec(439), vec(435),
        vec(431), vec(427), vec(423), vec(419), vec(416), vec(412), vec(408), vec(404),
        vec(401), vec(397), vec(393), vec(389), vec(386), vec(382), vec(378), vec(375),
        vec(371), vec(368), vec(364), vec(360), vec(357), vec(353), vec(350), vec(346),
        vec(343), vec(339), vec(336), vec(332), vec(329), vec(326), vec(322), vec(319),
        vec(315), vec(312), vec(309), vec(305), vec(302), vec(299), vec(296), vec(292),
        vec(289), vec(286), vec(283), vec(280), vec(276), vec(273), vec(270), vec(267),
        vec(264), vec(261), vec(258), vec(255), vec(252), vec(249), vec(246), vec(243),
        vec(240), vec(237), vec(234), vec(231), vec(228), vec(225), vec(222), vec(220),
        vec(217), vec(214), vec(211), vec(208), vec(206), vec(203), vec(200), vec(197),
        vec(195), vec(192), vec(189), vec(187), vec(184), vec(182), vec(179), vec(176),
        vec(174), vec(171), vec(169), vec(166), vec(164), vec(161), vec(159), vec(157),
        vec(154), vec(152), vec(149), vec(147), vec(145), vec(142), vec(140), vec(138),
        vec(136), vec(133), vec(131), vec(129), vec(127), vec(125), vec(122), vec(120),
        vec(118), vec(116), vec(114), vec(112), vec(110), vec(108), vec(106), vec(104),
        vec(102), vec(100), vec(98), vec(96), vec(94), vec(92), vec(91), vec(89),
        vec(87), vec(85), vec(83), vec(82), vec(80), vec(78), vec(76), vec(75),
        vec(73), vec(71), vec(70), vec(68), vec(66), vec(65), vec(63), vec(62),
        vec(60), vec(59), vec(57), vec(56), vec(54), vec(53), vec(52), vec(50),
        vec(49), vec(47), vec(46), vec(45), vec(43), vec(42), vec(41), vec(40),
        vec(38), vec(37), vec(36), vec(35), vec(34), vec(33), vec(32), vec(30),
        vec(29), vec(28), vec(27), vec(26), vec(25), vec(24), vec(23), vec(22),
        vec(21), vec(21), vec(20), vec(19), vec(18), vec(17), vec(16), vec(16),
        vec(15), vec(14), vec(13), vec(13), vec(12), vec(11), vec(11), vec(10),
        vec(9), vec(9), vec(8), vec(8), vec(7), vec(7), vec(6), vec(6),
        vec(5), vec(5), vec(4), vec(4), vec(4), vec(3), vec(3), vec(3),
        vec(2), vec(2), vec(2), vec(1), vec(1), vec(1), vec(1), vec(1),
        vec(1), vec(0), vec(0), vec(0), vec(0), vec(0), vec(0), vec(0),
        vec(0), vec(0), vec(0), vec(0), vec(0), vec(0), vec(0), vec(1),
        vec(1), vec(1), vec(1), vec(1), vec(2), vec(2), vec(2), vec(2),
        vec(3), vec(3), vec(3), vec(4), vec(4), vec(5), vec(5), vec(5),
        vec(6), vec(6), vec(7), vec(7), vec(8), vec(9), vec(9), vec(10),
        vec(10), vec(11), vec(12), vec(12), vec(13), vec(14), vec(14), vec(15),
        vec(16), vec(17), vec(18), vec(18), vec(19), vec(20), vec(21), vec(22),
        vec(23), vec(24), vec(25), vec(26), vec(27), vec(28), vec(29), vec(30),
        vec(31), vec(32), vec(33), vec(34), vec(35), vec(37), vec(38), vec(39),
        vec(40), vec(42), vec(43), vec(44), vec(45), vec(47), vec(48), vec(49),
        vec(51), vec(52), vec(54), vec(55), vec(57), vec(58), vec(60), vec(61),
        vec(63), vec(64), vec(66), vec(67), vec(69), vec(71), vec(72), vec(74),
        vec(76), vec(77), vec(79), vec(81), vec(82), vec(84), vec(86), vec(88),
        vec(90), vec(91), vec(93), vec(95), vec(97), vec(99), vec(101), vec(103),
        vec(105), vec(107), vec(109), vec(111), vec(113), vec(115), vec(117), vec(119),
        vec(121), vec(124), vec(126), vec(128), vec(130), vec(132), vec(135), vec(137),
        vec(139), vec(141), vec(144), vec(146), vec(148), vec(151), vec(153), vec(155),
        vec(158), vec(160), vec(163), vec(165), vec(168), vec(170), vec(173), vec(175),
        vec(178), vec(180), vec(183), vec(186), vec(188), vec(191), vec(193), vec(196),
        vec(199), vec(202), vec(204), vec(207), vec(210), vec(213), vec(215), vec(218),
        vec(221), vec(224), vec(227), vec(230), vec(232), vec(235), vec(238), vec(241),
        vec(244), vec(247), vec(250), vec(253), vec(256), vec(259), vec(262), vec(265),
        vec(269), vec(272), vec(275), vec(278), vec(281), vec(284), vec(288), vec(291),
        vec(294), vec(297), vec(301), vec(304), vec(307), vec(310), vec(314), vec(317),
        vec(320), vec(324), vec(327), vec(331), vec(334), vec(338), vec(341), vec(345),
        vec(348), vec(352), vec(355), vec(359), vec(362), vec(366), vec(369), vec(373),
        vec(377), vec(380), vec(384), vec(388), vec(391), vec(395), vec(399), vec(402),
        vec(406), vec(410), vec(414), vec(417), vec(421), vec(425), vec(429), vec(433),
        vec(437), vec(441), vec(444), vec(448), vec(452), vec(456), vec(460), vec(464),
        vec(468), vec(472), vec(476), vec(480), vec(484), vec(488), vec(492), vec(497),
        vec(501), vec(505), vec(509), vec(513), vec(517), vec(521), vec(526), vec(530),
        vec(534), vec(538), vec(543), vec(547), vec(551), vec(555), vec(560), vec(564),
        vec(568), vec(573), vec(577), vec(581), vec(586), vec(590), vec(595), vec(599),
        vec(604), vec(608), vec(613), vec(617), vec(622), vec(626), vec(631), vec(635),
        vec(640), vec(644), vec(649), vec(653), vec(658), vec(663), vec(667), vec(672),
        vec(677), vec(681), vec(686), vec(691), vec(695), vec(700), vec(705), vec(710),
        vec(714), vec(719), vec(724), vec(729), vec(734), vec(738), vec(743), vec(748),
        vec(753), vec(758), vec(763), vec(768), vec(772), vec(777), vec(782), vec(787),
        vec(792), vec(797), vec(802), vec(807), vec(812), vec(817), vec(822), vec(827),
        vec(832), vec(837), vec(842), vec(848), vec(853), vec(858), vec(863), vec(868),
        vec(873), vec(878), vec(883), vec(889), vec(894), vec(899), vec(904), vec(909),
        vec(915), vec(920), vec(925), vec(930), vec(936), vec(941), vec(946), vec(952),
        vec(957), vec(962), vec(968), vec(973), vec(978), vec(984), vec(989), vec(994),
        vec(1000), vec(1005), vec(1011), vec(1016), vec(1021), vec(1027), vec(1032), vec(1038),
        vec(1043), vec(1049), vec(1054), vec(1060), vec(1065), vec(1071), vec(1076), vec(1082),
        vec(1087), vec(1093), vec(1099), vec(1104), vec(1110), vec(1115), vec(1121), vec(1127),
        vec(1132), vec(1138), vec(1143), vec(1149), vec(1155), vec(1160), vec(1166), vec(1172),
        vec(1177), vec(1183), vec(1189), vec(1194), vec(1200), vec(1206), vec(1212), vec(1217),
        vec(1223), vec(1229), vec(1235), vec(1240), vec(1246), vec(1252), vec(1258), vec(1264),
        vec(1269), vec(1275), vec(1281), vec(1287), vec(1293), vec(1299), vec(1304), vec(1310),
        vec(1316), vec(1322), vec(1328), vec(1334), vec(1340), vec(1346), vec(1351), vec(1357),
        vec(1363), vec(1369), vec(1375), vec(1381), vec(1387), vec(1393), vec(1399), vec(1405),
        vec(1411), vec(1417), vec(1423), vec(1429), vec(1435), vec(1441), vec(1447), vec(1453),
        vec(1459), vec(1465), vec(1471), vec(1477), vec(1483), vec(1489), vec(1495), vec(1501),
        vec(1507), vec(1513), vec(1519), vec(1525), vec(1531), vec(1538), vec(1544), vec(1550),
        vec(1556), vec(1562), vec(1568), vec(1574), vec(1580), vec(1586), vec(1593), vec(1599),
        vec(1605), vec(1611), vec(1617), vec(1623), vec(1629), vec(1636), vec(1642), vec(1648),
        vec(1654), vec(1660), vec(1666), vec(1673), vec(1679), vec(1685), vec(1691), vec(1697),
        vec(1703), vec(1710), vec(1716), vec(1722), vec(1728), vec(1734), vec(1741), vec(1747),
        vec(1753), vec(1759), vec(1766), vec(1772), vec(1778), vec(1784), vec(1791), vec(1797),
        vec(1803), vec(1809), vec(1815), vec(1822), vec(1828), vec(1834), vec(1840), vec(1847),
        vec(1853), vec(1859), vec(1865), vec(1872), vec(1878), vec(1884), vec(1891), vec(1897),
        vec(1903), vec(1909), vec(1916), vec(1922), vec(1928), vec(1934), vec(1941), vec(1947),
        vec(1953), vec(1960), vec(1966), vec(1972), vec(1978), vec(1985), vec(1991), vec(1997),
        vec(2004), vec(2010), vec(2016), vec(2022), vec(2029), vec(2035), vec(2041), vec(2047)
    );

end package sin_1T_2048s_12b_pkg;

package body sin_1T_2048s_12b_pkg is

    function vec(value : integer) return std_logic_vector is
    begin
        return std_logic_vector(to_unsigned(value, 12));
    end function vec;

end package body sin_1T_2048s_12b_pkg;
